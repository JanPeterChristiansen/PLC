XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��2'E��8�oV��[��mw��!*��cO�lD3ޭ��0iy�^԰��f��.�B���4j=�7�F1e�����9$A�J�/ݴ�=I��� ��6����-�[�ۛ������H5M(&��}d7��Y���5,��4������6yH�� �X��J)ei�I�ϝ�X#5�sv�%.�����ԌpmC~j٭��<!S�D�0*��[��j� �hZ�q�Y�:�@���	�[��]�*l���Xl_}�XǘF������s�R%�H�v���c������4�\>E�4?ïl���J�vjE�����i<�EfnE#˖B�FG|����|W
��"�AK�l�͋~�����֩X�m)m�f
6��5<�{�q�/�xH��S�X]DE��Pc�U��g�a~7�s��B/HA�?ڼOm.Ū9Ŏ��
y��|R,IK�5�B�@+ 
����Y��i�{sB��y��~V�LǞ����Sc�EBP�����c�Z�*3���������zm�p�B鬱�{��(��3�.���U�U�N��I��A�`���C��\����:�����dXl9g�[�������%�Fb)�ȗ����m�|�v-s��³t�ڥlr�m~逢Ya�T��^��H9�E�Lzu�����J�� ~H�E;%9S��f����`7��{+�<���;���WiLp�XY�9f�@��&���{쟍���+�@�����NR��M�XlxVHYEB    c763    26003�{�l�y=$9�r�(�H�O֨^g����5�r����g�H�����7���D�˚N9B}7�������.��)��z���)G�%�	Ф��0Z�F
�=R�7��`X���N0�s�%+td'2sqx3����K���߁��Zb����1z@�W�
��3�j�b�u�P&��Ӵr�7J�7���0���f�T%�"D�@�X��ɉ!XK����T�qvbl��t6c���G�[���(��&�,DA�Ѡ��:�f��%�N� �B|z��{���ܭ�����IǀW8_���N^���8�K^ވ�x!n�N��`|D%r�m�`���2��8���Ke�*X�`[~��x.�T��|�A�Ҭ���3�z�.�4�B��<:ώ,vڣ�k�:��(&��1��X�T$ykº�oN%;YM�hi=:�.��g�Џ��0.�z��-�R�Τ+4�0�Hc�%���_(2��P�(�;=��=�S��r��W���`'�W5`�k���5Y����W{�0��sWc����؀��y��4�%��V�_e�,M!Չ�_ܕm<�0e{k��P���U��lVC��/U�^�㪢�U
�Y��C���7�g�gy<����-H�^fH�.�ܮ���nS�+yhY*���W���GAD�Qǃc�6A�k�
���|-�t���:X�����L�.�g�i`7������)}\�c����%���+(���s��j��<���b���?j!�S\E����%�1>�FK�.�Ns۰c�F��I0vS�W��μ4�;ԩ�}'��=G�m�G=�%���H����Jo�����'< s߻L�2D������_�G���ol���5�6��3c������� �X���{V��ȯ
����<��7�j�7�-6�U0�E��sYDk�	6/����'�!��^۳z�B�����_�q��`�%�oD,���8���Y�<��KA��f!������>:|(_��AnK*�� 6T�l<h��v?֝�$v��aj�q=<�̰%��X~�|Byt��n3g����E�p�ѥ�z��dؿ�g٪v��f��V�vQ׉q0���}�
����|�<-37J�,6�rR�Z��}�#�M&�_<m�0Q�2�r�X?U:к���X��to��)A������������r��t HK՜>�E�*��z]#���I��D�ƲF�P��8g��WN��<�q��q?A�ɵ�D2[�2d�d�Lzp0�
�q!�t"��/����N�2��PM�{�nc7���Ǎ�N�~0�ݳ��-ؼ&����E��ѓ�B*����v�lO�gdA܅����f����>w�v~���+,�u�82�8t�+����}��08�
�la��E�s�a�U�\?����A����a~��+��e1��~F�w!��可M�n�0,+����y6EaF�v�]��޶�� &c�N_CK9}�q����L��W��� C,v49�&�p<}���/)���=��*��mcMq�SΌ�ٓ�b��s�j#�Y�}�."&ĕ����J��Y,��C�yc��K��k�/�}�u�����0�cd������h�
I�HD�I��:Q���$�'*S]�mLl#�/��i�ߋª1�����9�&�L��\�8�Z��B�5�o�C��U���U^c����%��a�R7��)��߀��� ����QG��#�O������qEXw̐�#�
ނ���Úa����^�^�fZ�d�D��>���F�?����\1s��hG��I���ص���D�@3ھt�u�V2�6=F�Uq��4���6J�:�\�O��j�H�UȘ�Ί?x���;��l7������72ë�*s��v_�1�m3�(f2E.Ҋ�	.�-�0�tJK.)�fD�%��3�/MM�k���]y�~H�}~����L�)Nw�hB��`��¹Vkє1i@��F�'�%�L?d����O?�Uq�e����?jU�=��~B(�^���R��fhZ�A*�4ngJ��v��#�V���~^m�7�X�v�Mo�W�s�yt�ȼBp>�<n�ʅI_��!V�e��KKr����"u�X#�U�^�G��^a>�&�gd�_��� 
�u��
q�Y��-��*J%��8ؓ�-�>��㏳7b5f>1�<0AG�k��>��e�B] <�⏂!Q�{S�E�5�α~�;=U<��)�n����7��� `�� �E,[t~`�V��-����ĳ�^|��� UL=j������N3���GYP-�ϥ�q.Y��8�i>��u�!ؘm�	Λ��wC;���.J"l�����ꢎ|i
��J�<3?�3��b���O�I���p�s��ù_~cY�bp��p�4�����5��s�����b��>"DĹ�Ԡ{��'�d������UVK%b�ՎV���«�U�dXƃy�a$s}'*�<�9�|i�i�a�V �W���e);�j �/1���v��<�yw����]u�ǎ�W�H�!�*}&�PF| ���Z���q�;��#�Ez���yqr�6ZL�Yk�t?jG�[���/H�}�?�-r\����.���0��:�Ԙ�)�(��~�A���xk��p�H<�pd1��b'�ll#` O8�����we��	���b��Jy���)�Օ�EwD�5� y�]]-&���n�J�{��^5�p;�D���@��x��Rv�U��ϼӪ<)"�~��}��¾�>Y1,�������/�h@!
�h(z,�'NY׀�:̫H���d�@��ҥ���)7k��Q�p�=."q�7Ƌ�{+e����L�~D����O�[�NZ
��<-q��R���w�k�a�	��!�-�<�Ƒ4����7Nge��=<��7� �/�5�J��pW��=vsqEM��}�2V=B�F�db2z�~rT��b��X��� ��HIiT�M9.��<�	���k`����Q���b�o3���|6AN8C	��y�G�%�8��uKq̗�l����cE�S����Ɠ	�[�jo�t��ے�o�l�T���V����)��
��&���`�;�3A�M��w��S.���+G�W�`�^MQ��Z{:#�Z��>�]k�.���� ���F��r�{cRR�<JGF۾��a�#$������D.ul]JI�Wo�i�1Jf������iX��>�����կ����3�/ފ�_u��G����9��c��a�/M�T�!Y�JJ��^A�׶ⴾ��,?����"8�֜�0�l�eV�xt�5�]�'S��~p.��&�`��Ȓ��S�{R��U3��[�NH$6gi��1��\n��卒B�~aA����U��G*��;�4�:#K6;c: h����7�dNc�)�2?/�'^Xؑp��\��� �P e���� �)����g��hc�1D,F�9�m��\����4�2]0%�(�&b( ����d�ޤ�#~ժ��7��J�/}QS(�m|͜��Ɩ�k\z�w��;Yޗӽ�2Rĸ����R����%�q��,��8n���T��@�s@2�
�Fe�1��
J�5Q����_Z���n����8kP�����,��-5���4��cD!U����/ӷ$][EI$���/;T�W�_H6#�J�y":V'y����g��/`7���e���ٳVm*;�(�1ö�pPdQ�š}d�R�≺Ʀ�b\7lQ��J�^��7K�V9-c����0�W2b�.8Ũ�7�Utp��c��0��K��W`6O�x��p�Hq�Qh�I����!��P���tZ�;��d��b]�����Ԛ�}1��f"���E�ϱ\��aq����%+���y��k�i%��uW��_�@Ki��:Ƿ߭P̬#NB8Y"�K=O&�� ���"e�~�V�6;��U3�&�D����n���	$�i�Lk�"��r���]r��l�a>�'�ѿA�lѼ!��բ^�Ձ�NJ�_*�re�Z�Ir�Dit`vׯ\��
�;^*�g�kZW+�iu��#���+ad��m��cPEͱ�v��q5x��0u�\�_�â8(?x�B�K����������a�7�&Q��#Hk��)+�EA������p��i�4@C��H6�f[ʙ���K]���u����J�	35��7]qޜ�v�r�]�z��n��؛�"h�J����>e=��2N�~�`3'(����m�ത:
V�4s��3$�T	�3uw�d�D@0W�)�>�JjX'ɨ9���K���3�ǡ�MxoT̫��\����*[��|���a���7{KUE�$�C׈>���݆�!Ȱ���h��%���j3u\�%ًX��E��n0��;�$@�́o��;�m#5���
0w�;Y�e��g�����d@���bPyl��8�����ܐ���#߲!.���y�0$w��w�j��?�%��s0y����zlL��E]5-U���ご �eǉ�K�@V�G���4���w���J�D+�Dk#��ȩw���m�`ü/r0��N#�鯀Q�Wp�˯w��tq|�?U�Iv�&�^�G������&��K������Y�z�h]˥'A���$�{�BbO�4)��4F4�=���o:@)��;Ee�0�h&f��O3�<��O�b�5i�k7C7pnd�%��
 R�V��CG�EOCP��-�̻��lf�lu���<�,��M(�
{qJ��8^�;�����E�I�T��o�ɥ>{��8Z$����?êeM�w�O�@�9g�$5����F8��3���ie�E]����R6a!��!�{J,�~+�m/��}L'����m!?#��eP\�rPp��&+����l*Zl���#d��]��`El>��3%}�NF�vxQ�a�	]�x�J��ܲ��Fó�!��#�ϐ�����?��}0E;N��+q>�>�@�Q
�5¹Oh+���0p������L����L�Z\�U�A����s������RQ�6v�;��.��(�I=K��ұi[^�x!�����e��n6N�3��^z�UUI��{@$��7e���ݰ�D�-j�
�tiG�d��������lq����캭��ٲ�����1t��Pc�&��
��L��a�Jʾͮ��Fm��(��?v{韮���JJ���/��90��Q`�<�0s���<Jk���͸7�W%3�M��n�޺�0C��ŻՔwA5(e,(�CBu\yJjK��5>��&��$'CHnG%�U+��"��f��L�,z;���j'qET�U�?Dɿ��7yH�͡n��GP���'o�TxB��Q�(�`\�kf�S�r=�b�"���nMMp���Y���T�5M?�O^9��fQ�ʎ��8�j�q�]x�P���6��M�;3!U��q$����w�~�- 9�#bít8�g�BT���V��8��8�P�U�^�D�N�E	��{�pz�W�_�"Lt�8@~��dAD�im+;2�t��ku8<�=�4��q����f�	�H�!��_mU��KJ$f]V�5�r�x{bF����v{��J�'�d{T�������Ȗ��PbfP�� �s8xB�ە=;���
�{��(�"='�����a�����Ԙxj�9�DXD� �W�D8gX�{S^B�&�T[=+k�	m�����r;�!�a�'�fmX@��@��]��H�IЊĝxM����>0�Xf|�-İ�W'	�B��Ί+�G��D�XX� .L�Z�y��fT��| �r˞�A���*��w�#�K2�F�����=;��y�ӡY`a����#A
�	��W��\ƥ��xZH�d"N�	�</fy��Fk�[j%{��Yc�An�Z\�,��1�T����*�p��L���ރ��bџ�a�0&�φ�G)`
���8�Ҍ�׮��=��=��M�1����*���,��Y�im?�� �̮o����^��/0�q!8���-�Nx��&�$����0��/4��o��V�_Q5нq��1��, ��Z�`��ئ��5���d���d���3dD��E�����p��f�N��$�Q9�{�v�� `���v��D�O������.�o_0�{�^5$��U�7`��<[#(�\�t��:^� Yc�������8�]ng]9,�r�W��\\Ed&�p�a�Ø8m��A��,���JT��DT����@9f���"�$��C��ۤI0%E�J}���|=����-�j�P����;�~�?��x��z��tH��D�w1M|9d�ƽ�佭^T$���RO'�}�6E!��Df��X�@||�$@�%.�� \� WZ�O�U0�]��u�sI�>3�؇RJ5m*����G9���E�>ԽI�hS�t���^X���<�.'��];��(�E�_;�C�o��aq������pNl89��ݮ�v��L�����M�����:l�h�
�i u���s�暴)~[udC�ၚ���ƹ�3�4��d�*4T�k����P��hr�X�ݚ�]���tm�Y	k���Qو�� F$z61��ش�藫�
��^r��ş�[j'�j���v�"��	�D�7K�(��-�#�:�4����i���IGBQ;eS�Ϡ�P۽��X=[��[[�|����+�8@��0P"���W��i[6���_����0uQ��!��2%���C���[~ÂO����R��+�F��Ry���X�s��N�-CRYX���2����΍]j��XO`D0T��
t(d���~�/u�)wu"0��tQ�|֔�HW��Qp|��D	�v��vY�k���g02��W9���9��Y&�Nԋ�I�t��R~n��<���a�}�_U���l_�c<�5�]�����<�^f�>Nr����"�O�'S��9�t�EcS�����P���h�*C%���)@E��N��t�

+�n�2�eG�9 b������ϘE�,fx��egv��>�=oe�)����}
�a�G5���Ќ�r�8<� eA��S�����듮�O����d�)��ySי��b��Q.|��
HEτ�s8�ԍ[�b�A��s����zv�|�A,֙�4�h��ホ�)8�"b����#�jL��`oɥ�4�,��#�m��Dx�Z�E�vJ+�'�5�W�(<O34}�|�E��l���*���xn}b$�W�@��#>s���VF0�T�(�L\'�M*�R<,�����9�ሕO�A��a|i%�r��w��We��_R�D�ʊTI�Q��CDU<|���.PiО���qJ?��
�v�F��Ҡ��]�!�����O���?QS�nɮ+t�f$uD�9~��o�w����B�krb�v,*�l)jsGC7�'����(��q4��{o�e��Dv���U�^`��R�I$j��@��0S��!PH�߶2�bJ)�$���y�7���+%���/2IF��*���¸1���2��Y��v�x��c�S
J�`q����[H�l�gL߁���ǳD�K�ػ[h�+�է�k0�D_�N��`��u֪I����h��ƚ��=8�XXR��ȤeA���q]��m<8ڠN%����Ϡ�	)Y�/�����U!̛<`�mP@�E{����Ɨ�c;�d���{^���V;Y
� ��=�Щ`�B3iv7*��T)%����q�|�
����!��<8�6��%�FX\�M�	������?cǸV9�}q�)
�>,n�ٰ`k9���*�zɯ�}��(b��E��I]c�SdF`�Od�BnOQh=�-ٔJ�����i��q��v_�������fsi@QӾ^���L�Ҕ�^G7"]�C+�2� ����ט�<����N�T�^�ޅZ�L�����>�#SYZ�+?=0a�D�bF�؉�8�}����Jz}��j�B��"���Aԃ"�͸o.$[��w4��ƅ�$�?~�[Gp��"���Q{jX�j��7�2�C��,�d|��Cs�h�TŢ�Zv�������JD��LAv�KgR�-u��evE"5oF��W�4�6n���b+��ګ8��;���QCg@�sIC%�2�^�<M�y��9�%A �Y~]���,����*��?o�R������ \���)t���{�1�a?�eR��5ٓ�|�-��즞��� & �#�b `�&�g�!$�V�c��qT�.�=�C�S���A*�fm�..|?�"_hk�ũz{,ԥj����gޖ u��EXV"�w?�DDB��t�I�	�v��\��*�%��4�ք�(:��G|��pnf^�rA9=�C�(���FP�TtY��擇U*{g�Q~�h�d�`gxbQ����~����O����S]�L-�~��I/j�~[�mV�|%c�rC������-��1`�: ����R4����ulmF/]%�n̫\���?�. ����y��7@�:�J�RA��0�����K1��$��1�
׻��e�i��{�HQ.n-�}�	m�u`'�HS�s����_�96���Aʸ=F_���I�cR��'�����L�Js����@��ޫ;���l/;���@�q��*���zVʨ��b﹣�4�W
ݲ�;İ�"���(����w�m�c*���v~
�4� �u*e�/����0�����{۹@%8��c$0ñE��`�#�;���M�J;T�:ۑ�m����3��0���[⺶�M�#�$Iߐ��]s�w��a�q����� 2h��Z�ZtFq����A˟�%+�~�S��a�p(ݳ}�Uuvme��Y"�H�o/�����>�:x�-��V����y�6D���ۓ[+�*��r�thf���r�5��X�:7.]QN|��~��f�ϊhs���	S� {t���grۘ���4�j��{��U�Y#X��gH��Գ��')7ny��|6bᕠ�Z���ޒ�Y������>���~�ȳ��E��i�,��ept��e	FK�������IO@7�~�頚���-��k_9�T��C�h~w��!��I���mJ��M��<�3$�C])��<�4i����EJ�2=҈:~�ۜ�������x���09�=h� ?l�C�|������Z2s�f[AN.�AT{�.�a셯��m�i����R=<�~���e6�,���5{�=P�ȫ�����ͦ+0f�!܆E��vs&̞�)��8cԒ�׽Kq'�5w1n�Q�d��Jҫu����h�	"r����[(��CM?���"""L��<b�STB�<2���ov#�"����3�X?v��DOK#[=s���8��C�&���dv�M����t�{Wm��~�ro��J�b�{R}V���`��l0u�r�m]@���c�}�J}���n��_���=Kۇ�!Z��f!R���B���w?����m��A�a!�D7oGi�<�PI!]���Y���f�<*�Ƅ���W#[�����	!Єlk5g�y����)TF�0����ۭ
������I�ҩ]>t�B��&�]��Nj�1��-�s�(k-��;d�
,��ՠALҹ�ǧ����0�B��U�hq��]�"��͚T��9�sc�S�A��ڵ�G���5������B-(1B��G�/�T�����Us�Q_�o���Qi�Y�:$��T,�w�ܒ