XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������3�]ӑR� �B!up�Ŵ���-�+�����A�WP��t��)��Ck��P-i?h�A�N�h��ռ�d���������K��JtH=jAB�������8DQ-�?~�S�	�?5(��0���g&�9�:�ͧʝX�i��WA��+��5��FX�&tq�.����C���i�,`^�Q�P�2#�6��^ ̮�����9]�N�Q~���|�9Sm|���3�9�8$_t�	Ey��B��މ�<���Fp�/VK��fT%Pϥ&&��BR �-MܝZ9r\�&��t�6�*���u��k��}1D��'��.�����4��0���I!��ܯ��vܹ2Bi����ߏ���ofcJi��X5�$�^ �d�zs;l����q�	SJ rXS�dqYr�@�HLB6O.���=�C��g�?���@�F�*=?��3<������o���������sEBĤ$�փ�T��1�ʼ)l���V��Z����6$}i�[�<�	�yq���s$��N�������Nt
ݍ�*
o���v�@9�i�9:ʾt+ݧ�3p�.E��"Fo2��f�	���	���:�"�~�d�9�A��/m���T���z����#��@�hF9�&��p�ow,b`��+�\�]��Ip�I��Z�j��2o`�B2 � ��*�&�������bes�Y�6J��1����D6�8&�\�ҩ�|&�B��v�<F�ko���[�0X'M��_�E�/f��<1c�8��B��u>F���r�:�~XlxVHYEB    fa00    2260�=��٦S�iwV����F�<��c�
�Iq�o��!<Mz��x,����L��]@.s���Z��5]���&,��S��yz���gjh��~ub�Ю�Vϸ�Z�����J������2Տ]`��3��^\�rV�K�K�pû�X���<�<����=���7t;r������Da�Ԁ�C��8�]O$��T#r�N���ŷ$<t�.�_�X��P\��o�w�ԏ��7��A}��r�%��&�L!���vی��>�!�-��n�&�c��~�C[��ߋ�>�Lo��U8ii�bz6�sE��WIRRr���}
�o��K}�c��*����y�,;�^-[A�B��u���J��mŜ㡻<	��Ji��z�����>G�pފKϏ�^�X�6�>�.�������;R���.�U9%q�������cC����B���^�����.{��L)�����k��N>�{����pp
g�#�w���׶���{��vr!w^loz�V��HI�%MZ�ZT��封�-�<�dU!�OXe��Dt-�N�E�^)٫��ݣ��0��
g3��l2��@�Pڦ_�D�_f�y�z�"���<�iaF�	�������$6����9��#E���޼�9��)�T�N�mw9tF�ʰ��B%,ީ���&'shL�K� �/ ���P}Y{w�x�X.�G���6�5�j]PFΉ8?�T�2j1�E�2]6��c<t�������+�p���[���=�!��U��?�b���1֊�\O��,~��cC��2�0���Y�M�>;)Ȳ`{=���m�L�1���:F|�6$��d�Ķa�D�t�@lfq�'��
�L�������B3��t���y��7J��
�Vڷ.>_���|����5�=��X�BL)��q|l�M����{�(*�;�ձ��wC�i\x�>�63�!�>�S���rY���4gi�o{h�G��㘱��L.5mY�%�:%�H���F���VX�K������G��06ivvt/�#'I}C��61�>���ǏR���m?,\������t�Y�R���;e ��L\�57Nx^P��C��#��_���Ǵ�ԡ<xnTE*�,O�aJ.�lh�v'�8;w�t� ÂC�ፅ����5�F�w�گY�~��=��*Y-�����Bp���o�ܒ��n��$��N��&�pۈ��H/D	n�%��֪�8�{ӘlDwO�P��&I4�q����ɫ�WH�1���:u�y_��R4%;���e��BK]@1@	2�W�[)�w��;���e,��3��F.0C�]/�Ǟ^0�[�	/�QZ'�������(�.n����E��V(�^b!�h�;��S�c��O�hf�����#��(�#����.(k/Z�V>*�'����vz��|�	r��:��_AW$�Nz��z�/��9V`)m?C}8������_v����� �\'Ux�ʢ��(vK���W/�E�8��g+ ^�y�o�iD6�e΍��,K�*{Qs�o��ؒE��������#����K�
� �ݡ_1_�Z�8hM�LD�fnj��#�ϋ2Z���GV1B���-�F�0)	�7�y�J�E�C�\Q�{��*�r)y�@ݭ�^�mZn���'���͸�˙�d�<P]�p�HD�6�3M�ϋ�j�gZ�C{k��&�X��}����xUW�s��
~�vL���Z&^�7��!K}0ṃ`f�d�T��:��bݩB��e��_3H�OY�I(�uO�P��J�/�oi����_�4=�W�j �B�<����DO���It�Iз��d���ol�S�4⁕/���/��"�/���Y4�L��T�8���y7"$�~Z<���'UB���2$��޽VI�k�!Fc�m�n���N$��}]���&�$�<2��?_��ҭ�e{�,qn:���7�Z��VK��9����m�5�ޘ������0�����_ΐ)u��H�A.������|�#�`ޱ*�V�"���腛wɩf���FZ���z�w���q_z�|9PҎㅃ@LsL����%���U�L����#�T,1�F60U����sS߂}5�k���|���.Yؖ\Y�5ؚ��v���~P9*J���.u� �<�6��<�E�!)����`��[,��D|�G찭ݥg8�KtG�.�-�֒߸9>��s�>����s0�im���GE��ԾoD��̆!9�S����Z@���$��'��+�K���j}pH��!Y���_�шx~��aF����"�''�w���"0οcU�P&�=�d~�c��.�{�n�"9�����0�?.��S|7�c}ƈ�_(�E�58��{gT�}�H��OdM(�����I51�칫��W�-+�]�����Tn�a���z+����|��.fC���/,�M��f����je}m����S�o�+A�g#vda���]�K`_�X�a��p��ф���%b���*��x=	4ē�����i�v�ܦ�=�2����7z�
�7+�C{?�R��R�p�sf�ԙ�3��*�+��B���|�)��f(�߭������~�y	̓�J�|#��r�4mCy���C$�P7@�_����;�e@W�l0W�Pe*'cNKds�e#}<Îz٤{�
����Y�l^�0\���XT����ϯ��4��.5�^��$�P�UTR^�\G?���P����4F�J	w���>���b�e����&�:����xԕ $ӴL�|Ћ֝	��a��VV�NJ��X"=�<_�Q84��)��x!m����Bq7 �� ����ZR|i���E����S��S,��p�Nuu o)mv���^w��U��ŝ[�b��>��W}źI�VK1�_W,nJ�V������+T�����LP6�Pe���4��6��+��O��G��	��S��Y˕q���[�ۅJ�f��K�S<�d �]��!�/F���1�c^�Ի �s��x��V��b�<&��Q<{�֌�u����% *�hcG��#I�d�sjk$����o��k��qG��Pq�W��Y�n���7��X#vx���k@����ѐ�4 �����/Yk�},S�{B�'
�v�dI �d�l?2E_��]Ge)w���7U$q��MKQ�L��e�6��Ȭ������K7}(����w�	O��sΝ&vO�φ�4�m,dJ��#�[
{&�q�9�a*@/�j�+}%J����%�~��Of����=�'�X��vI@�ܗ��d�g�O|'*�W&d����w]2ИD`���<wT�/��#~���…���7od
ɭn�)��hɤ&�4���j�����\T��Otb����K�O J�L����Mr	���dp�i-�/X	�#x�*&p��L�9ʩ�����ZQ�ҧ<�ߑ�b����Xc�8gHK�klͱ�]�LKM|�^>↸'O��9ր�ϖ"�g�y�ߛeg���8� �S��� ��B����,�� �&����j�u������uW��S#^J��ρ���m��9�-?��S�Ȫ&��z�&e����<-���������|�v�r$�����,j�mcB̕��#R�o)��1���9�f�F��Q�}��?Z���m}0i+Y��s�Fk�4g܂��1�*-�"�ӆ���[4
�)9�]Z?���v+�|nu����K�"	T�[����U+���L��I��Gc����ɝ���?�x����C����)rb��WY�<��_E�k9w�jԤԚ�b��/؁�\j,QjXCU3M���ѿ�@r'C�����L�	� �/���o:���RE��e*�A���<v�&���3�@��U�(TZ��9�U8�m�ap��k��)�֭PT�j�~�<Jٝ���sr����F�j*q�绔Q�R)�uU�y�n����*~"_0���>R�^��B�x�����"��R�:2���Q4'"���ʸNcSV
,��s[�~�Aai��jĵo��сs]�Q��3��|����*��a�Vq�0;��J"1z���G9ß:��ۧ�W��ͱq��x I�+�����X���%\p�2F��~0��9�
�2�"�/����,�Pﵑ�vk�8vvO�g2��,04������]�K���u9����*%�W�F���E��h)�ٶJ<X�� �a�׌���i6����޾�"H�(�ڕ���i���@�'�Q�%?� à��f �@��?}5?��� �;���.��l����P	Z�����{�5�Y�ٗ^��4s��Q��y�ꤗ܇�}!��k=����n�=��<�G�V���`��u�
�3m1}Mr���h2�A�Δ�Ф�%3?D%8\�b �C0���th��23I~�L�^u���^��F;��#0#x�!d�!��ƮPw�8���o}X�)�@�[<q�;Za���1�[�y�l0З��V��7�'�{����^��5�=��!�tT�;��D�|���渘}�`������<Z���ԡ�H��Ja�ޔ*�>���ȴ.PҰxs9�tV��4��5�Ϗ�z�_9uqM���:I`F��<=��@�J�Ւ�37L��!�YhA�?W^�)ޞ��{>A0u�c �*9�MA~<`-�j��5�X*^���2Z&+c�,�Yj�	W�֔����J���S�m�q �-R�[�ꞗ�U���J	�/��&$��3B��Wc��n�A K-;@�9=zw�!��ː��Z���>/�����
�ԶO�ʇ�/��H�\� N��z�V��L��dNp�rF�T�Tm5J��ά^�wT�y	h��2J�r"� 1��-	������߇R�\'P�zT�uQ�\��\�E��(Y��W���C��4@��O�<Mp�XL(r*фh���Br���	+�wϼ��I���rԺm\�����V"W�HY�2�ΰ�l^���k��(8�L� �OVؼh]f���4��ػД\q�LՖ�g��x�c���U?*�ոw���c��� o��K#Z��8l���Y�י�-��*c��b�'�0%lEv��3ҀJ���߮���/p\�*u��z��~��˽���J�ۊ����� ��j�߾J
�M��ɵ�|�	�_��5��Q�Eu�"��5p9M(]r�R����Fq�[�6���q������i��M�U��#R(5xq�Z�S�/�f�T:�W\D���ɮ�^�\�C��~����i%{!j%x;fe�;q����Y:)>�����M6�1
�X�m�y�P�g���5S�d*CLx'���L�Ңl���'�B{1R�g�q�"���	*�Z��ty~H���M�ؗz��E�N.ߥ?ԙw����U�}�Fs�P_�t��:9����nZeY�;�+��B$ۨ�X5�Z9A3���LQ�S�:EG�.����]a���t\F��B��&8κK�N�m䦲��
�d "�r�B��lB����֖R��<v��"ǆj�@ӺQ����DȘ��(k�6�q�����(6DԀ�� �8ƨł5���?��d-��h)���{���Y.R_䫝��|N�Q<��ʇ�,ч�Tn��@�h��l��V��R��"���-�O�s���K�X~���DjQK��_frM�QN�<�uX�f#z�`m�so�E�LㄆBp�G�8c�{�0_��툯?��PZ��Ǐ)�^TfOM|+D;�3od�h���;IK�^P�V��m�z �Q?���C/�=ض��٧פ24(�Kr�L�>GQ�*�L8K$�yUaK��G�=�>�9�HԂk+�I�^�\ز�Ӹ��1�޹�)���$�I���[��.{k��\o�*B�v��j�Ԝ�dp�]�ԮFU'1��������.p7V%�������>���/n{���;�oi\p�ߡZKeb����9��,g�gg�����<�S-�hBEL=Jr+%ya�v���g@�'hn���Ӯ��ʍ�#���#>D��Q�狂�Y�֥!�Zc�Fpy����̵��I�kY�Uz��#���0^�K]?���0B�L���¨~$p��6I�<쫪�kj����D�6���O�'�l�۶ٺ)��R\K �����*z��9�D�_��!Ȍ8>%�3���A�F`/DA?NV����KN�u����F�ذ�	��y�!��E3���z�a"
DZz���U�`�������-�b�H���ͅ_1ґ��(�8M8��R�+������4���=��ش0���7�����U�F��thoi�?�Zn�l�/?5�� ���3�գ��c&���J&&tq̗	�G�ۉ �AV�V��y�6�|��$%����y	Lg��F���p�T�t����Pc�!�ӭ��M���;�۫��z^)����w � �e���P�����X�X$�l�c��敮I�CM�7wk��H���Q&
qg�..��$�K[E`o�� �N�ĈP$o;Yb(8A��>��2�g���;~��V�^��<�x~��n|+�, �v�����o�tX��+T�N6����òO�O2M";�ل�es2���:J��q2���\\un�A�}��� &�$��y�&ƞ˫N?�ޕ)W��f8lo�����-�n���*�_��E�+�>$�(�l��)U,��)�qt�Ίۡ�Z	���|墧��x����E ��˳�ه鑕.�[�1�Ќ2�ȱ�dX�{K�	M����ُ�f�
���������0�^�u�Y�P�^`Y�m_U~.����_��@% @�R�g�����w����F�S�~�1A��5�	er�|dF����V�J�+)#�l\�p6ꜝm[F{o6>�o6E�мy���_�%wq�{��c�n��M�Ū�G��仼�o8�]�����%�rb
��,�S2��W����,��ca�X��1�� e*�\Y\[p2��b���� �b7�L�,���{#�������qI�}�*���x�Ϻ�'��8����NU88W�2b_����0�sk����[�����m���R���U,wT0U�@���xC�E��;'���bt��*Bpm��>�s�έ�5V��?�oǄW�Fn?ɭ��S���ϰ��H�l�����[��tnw���)�=� T�߁F<���AR��X���!�DV(ہe�U.�E��x/�G2UD8����0������WaA�@-#<���D�i�/MV�����5��+yy&/H�&���ԁ:&�ˉ�M(��&�
��:I8D&z��P��M��ee͆q��b���i��L�c��V$�p53�h�b[���M��5y��ܮ�\��bz��\::?$�q�3����7�/��^[��� 
2����v>��h<�XY��cECaJC�$1�d ����UA i��9݌�F$��z�D@�8uh�A��K��c�	���ZjH�;ŀ��5�9ǫDT{ov��p������0�}7�����i��P�[D��%QH;vC��ة_�Px������pH�����l��x�{W'h�07�ʗ"�i�,�?溰&s�$����FZy���=��aN��	/z�`;Ş�6@�Sl�c�<R�kU�{7�8����Wi������bx�mǝE�œ��#-�����9|�;lj�-"���-���I�}�(~G�1fv����=�!����&�`�b0��ug���)��<;�n^��<��]�ڸ�W��-�c��b�,�SB���~�x�u�� (:�xl�L����0^� �e�&�1��<:!z�I��̸�܃�.k�@���>|oڇ	��1��d)L�6�C����~%~�J��}�I���Jn-QD�H�jt>��r/q*��VH	�"�����X���� ˑ��j��?��j
ήv�"e�n�,o-v0S��?��uQ;&?T��,�ُ ��%	��)Q���l"J���9b4�JW�z����H<��pu�8o{���O�y8���='�d�[�Μ��z��{�?�6{�:�r��Ŋ��wm!�C� d̑�Q�����7�-�J������T@i��L���j����A���Me*H��Ԙ|���r84}ֽr����QV�{�ؑ����09�GJU>kPY�,��#��L��"9��6�taH� Ix}�,��Uuf6Π�7����S����S��U�ZQb=�,8������Ꭰ��\ h��usg�!�5ʌ�#�"�� �v�]�y3~�B+������M�B�u)M�;�����`���Z�i���[�g�*��V�ʫ�^�״��>E�����$B'q\���4ڽ#U{8�Fو��n��ՕdD����1�/�\E�^j٦��~��ֲ-~G,��fG}k4����&5�u�$,g�F����W�.��h-��ͺ!�6����O���8�MT��Ta|b(`>�$�Տ�����f]_��%�$J�ð�*��e�6�}�A]���up>~p��N�z�iI��[Ue;�
lǳ�>h\��7a�oo�]��G������&�.- �����n�eo��Jq@�tfa�w���yu�℮�=����*���ѧ�>�ƬQ�|��gga�[Q�T�����2�;H�����[�UT��Cr9ԫk�YG�`	�
$g����U#}��H#���ja-Eس�N`�XlxVHYEB    674c     5c0�[�����2<�}k&�'�dZ,��Y����p�J��ϫbY�D�u5���<ݸ1*�x�o=hW�$h�6 �n��޷��΢#~���"�� �F�i����\��}V�0n��@::|<�aT�g7�E� AjQ#�7X�u�NXa�F�B�)��zk� p�b-�Ov� ��4Uįa��1���m��PF[�=���w��#_��6���N��+F|b���YL�8VɆH��c�i�	2�V>�(DW�b*�F���`]���9�_�ۻ���x� �e�@�i(/�M},L�M�ڳ:c9�����B���B%�S���V`�A*��N?�8� ��m>?�x9�uG�e��n�����dW���|���g���o
I����B�3��+� ���d�U�3y�[D�e��d� p�,L ����Ƶ�����|���ntt�-�3fv�g�ylԒ��"G��J��q�1�D-Ҹi��c��@W�X[�ODkUP=���z��'#m���u��rnI�Q�/
+e%�܌6�uڨ&f���Sj��F%��&���{E�&=�d8)
�V�� �z�[(��}�7Wc��Cz��?�)<����\����b�5�S�ع�� ��:�����Zw춖&g&*P�'��ZB�Z��R��C,m�5#�(._����q�� �t�#�ý���a|��o�BS�:�1��Y�F.��5�R��J�U|����YL ������l�{L� G�rq��b< 𗘸�c��\��������NZ���O/��ZTuDX���2$´M ����,�f��k���=�p+ƛ
�����o|��1�X�-(N��ж��췗����WIj1���~98u�-���#���I�SRl��݄�*��=���Sd�~% ��0&1n1 J�5p�J{�!z��bt=r��q���@/m���BÑ{���l5^pT��+�T�<.>)jM-��͠��Cf���ڧޒ���k��?��T$c�?�=k�W�S�n^�p��2��ؑ�	��C>ؘ+*������u�X7��7wO	�SG�C����qc�xR��*��������Y�a�R�H�ҡ��a�3[��Zɣ"�@���5>�/&y���)�>b�9N����l���B�lHdD��)y�F��R�~ț��PbT�S�bTJ�pR�0Jb'�<n-w��G�*�J!�
�m�C`�9�-��C\�����$��aX��8Mt>X�j�hn�y��ˢP�)�B���_,�w� qA�Ћ^��1zmμSuB�Q=S=Q9����y���2C��mרҟ��	�f�s+��|T<)�BnD��n���g:�2qo�����m��������|��j7ͱ(D ۨV3�͸d���_��Hۦ�g�i�D4����L�0����R2�&֕a{�M��}�M�6^�y������[
x�Ģ�s�������,��w����