XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��H�E,�1��E�Ʀlk|P�@������l�W�!	�_�:pK�0�2nEO(�������>�MA���M(���B`������ө'i3\�泥�.�yl��IpqK�\#j ���������v�~�w�`�W"jPzX�>+J���'�&���t�i��Gz(vH ��M��P���	.&��ِ6zI�]�#O��)�1QaǢBj��B
��g�r����6��)�x�1�*V_�r�^��2ak1��1:�={�el�Nf���!���B
���8���w�x���q�Dh�p0�-p����7Mhkھ�<r�T&  D����S��'� d��0�����S[{a8ƑI���Z���ԏ|rD�����r����/�#��mA���l=��.۱�7���_�������'�6đ;7=������3v)�8�oԃLR��x���/���ڶB�����Ŋ��g�:���1���JĎ+��pW�x��
���.�nt��y���n�L�җR�{.Zq,�᪀,�h�D����,X��6L�z/S��=���r�{���"���C�C?�.��9s��/��\�}�ŏ������#���\���V%A���P��kt�+�J.������>��Ӝ��J 0��.�n�1W*�uj�Sջ<6�K(��ȋC�|��:_�(K/�q1��lg�$ad���g� ��/���	��m� 2R��닆�����yN�����֠��!�OF�����z���.�XlxVHYEB    9de1    1670��@�|ٺ�ܲnCS��V�P�5mK�M�p�d���o�B�����\��c#��N֫����H�ǀ�PJ����-gYxt�`��Wbk*cT�j��3��a
��zW�f��X��]��H�{��SƧ���o	[��+n]+=��������a��p��C'�;0�dஉl�������� �&�1w農!u�JP�c$ ����8-��v9��,�,l�w���H�{
H��t�5x'd�x&�eL?O�&���'���E=\Kb�5�V5�`�0I�s&F1352`fY5د�P{0��*/Vh؏�y�����5��o��ȷi�ś��O���%�h[ij]��~��fG�~�J��Α�Y�������W�F?RS5����ӝ�	f��jY�r�6ֺ}�֥Ps0��g���i{�8�5\��I�@K���7���}��HY���Vb�$�E�����bB�]����PB���*���4��gjj�z3�a��К�9�M8	o.詸cTOI����ĿA͵�����0���sǷ�_���&Q������ciQ��}V��	���SuX�G5�q_4b�����r��t�c4¯��"��5�t�C_G���G`���y(���$�˛؉�P��KV��O�c+[c��WӉ}���pv�w�c����u5	��0�� /�E�ة�RO�&�C�C[rh7�+Fg��{�._��Wى5Z@��r6K\.�i������Z_I��@�+0,`�&�$[i~=�4Tu�eN!�����FL_R�`xt�����^
�f�/h)��vk�Z��l���N4�}okA�5�ޘ����{+Y����7����`�؏���l�3]�df���XO���J���G��E#���(k���a����5�j(9Z��M�.�mL" <��!�|��~�gjہ��������.�����X GG\ΧF���x_���`eGC�E�(�R�~�Z��0]��K�h���X�Wx��)��C���'��� �����G�������I�ԑrb��kI��i^�t;�+��d�.�*Ih<ǝ��޾�-��-#`� ��:��ʔ�I� �.-͵=t�>�t���-�5�/a0��Q-4�>���Ӷ����KHJ�:�vY��Z��X+
�3y���;	�E�B��	��h�����FN���"�>X�0*Rv}y6�IG���sf����n��zT�e=q@���4aiѨ$�Rj�uih�n��(k�� �V��R�m���Ʀ��\�*���˺05'Y�{���⿜�����]gw�a�XL7�ӈ\�<UO��F�.Vb�2W4V�G�d{k�w�;�G`��'`SD7CLΩ^��h&͹���Y)DE����N�oS ���ޝ�|�����-G=,iCo��?*G��g'�*���iD5g�̳7~��"h"�T;b�߯J���=�׾=�k���u3�x)��ې����G�-H̉�y�"������X��l"��@�G����m�r�� yԌKKhxJe��H�;�����?t~ ?� n�Ь�<?T4��'>k�_l��0�ߴ�$�� �����<�9�š�a�ت�#��~v ����6�]��+�/�Ah�V�r^�/D~(���4;��n���C��KP-vP�ߠ���'��&��/k,zNH?6g�>L��e�c
�t����p���T�`�C�:�{��sI��_p9���(5��h��?V\�y��e���%���{8^�xԋJ���1|���fgTl7�Ң$��z/����=��yx�dе���UQ�5Z3s^J����R]��Y&9�A��(��M���è��� 1j��;�%a����"_�Q���	��1�����3/� P���B~m����m۱~�b�G�Y��3Y Ǡ�hT�b$q�&�z�x��a�������!�d�tA� �1'�6v��+��zi�mp.4�6Vq�٭@�OL���<j�<@M�W�%� �����/���Q�!jA����z����rQ��ۇ7����".�qR|ۋ��إnJ�,*���_�\Gd���'�3&e��4t])�R���s����P�j��!l�B=��s'��&����2N�6�'(���;B6j�	��_2��nq��C"�,��AB"aT�����Qٖ��0��<8�I�,�?n���|�ﶫ�����Aͺ3���7#gou�</��&�|���H>��L�@ͯ�7�a}�ݯ�!��Ն(6��C���U�j��q��j��T��V�X���a]���SGC�f"��ᜅ�}=�L��㢷�|�gi�ߖΛ�l=U�Q�����9�R��I6���r�~x�Y:jwXʙeY��z�Y��[�X��)`ҳWJʄ��\�[���L�~J՛z�`�K]�x�͜n�C9��W�����e��w��
����3.Y�6�إ>:|iۗ�3����ꍽ��m�R�iyo:� ��y�X�|��'bA�>�.N��k�md	�-v;����v�BϬO�ú���N�l���/
�Ḩ��A�V.Dix���D��(�]3��F7:��veOr�@j~/ǫj��6�X�q��v�!G���(e��ooG�����a0q/CR���!��C�A���A������S��'�1*kA+�|T�},X�sH00��8�\!��y�w��G�@=q�����J��APY��~��l�k� ���߉a/��K����)�Xg��%�{�G��/V� �c1N� Q��:�_�Y��6egb�ؐ����G؂Cşl	�3���G��&z(Gw��׀P�h�-j��Z��i�z(��0���3�,b����X
��$�I�{D�#}!��~����e|�GF�G��Ψྱ�9����c��6�|<�M;y�s!�1�5,$�b4�<���]�Œ �W�P��v������8���D��DŘƁ��L��e˺m�1Lw��,ޢ�ns��^C�Z����D�4��*�?�}��pv��f�kE�U�	�ъ�/�%@��2�����e�s�=�$��x������M`j2DF�~5���ʮ���{骰����;��n|���;�Ŀg���![���a$���w�G����*�rv�.��])�H�M���6�lV�߶|5|����Ӝ���9�"#k�e��i�i�{Qw!��( P��%Jc�@��|n)^�A��%pXN�ٚ�3�j{��� ?ѐ{f��*�Y��}���{�h����U�dѩ�b��m��ωs�&N�ݖ�J�<aDN�D߸���^�K���N��=@C��Q*�f|S�מ�!�0x%g�;��7m8%1�/R6�o?K����W/ɢ5S͐ $�ı9��.6��f��m�Dw_�SHj�j|-q,њ�'%����h&SI���Z�����8�,$lc�v��݀|fZ��S#��p��K4TDg��ֹ��M�r����;�@�Ξ����)�}�����Fn�=D��S'H�5�4�ZJQ��(ݢAɺN�l�`���IĴ�>����^�M�Ky$��$ٹ,b�	�6�})MH���w����������ߒ٭����$�A׿״ aUAF�Z�M�� V̯sA�\Jf%�"UϘ�#�.aA�hLq"h��3���ȵK��p�~º9�ز���b��O$7ڪh�X	5�3jhf��Lߥ�h��q" ��L��}�/��w��pF��s}������.�pc>`���r"1&��ٳt/V�ZF���p��fW>�)h����?w������H�n_��ӛ��������0�zF�o��CǺ�
���}̅@��q��Zۓ���D��4�����ވ'�xc6�R
�~��#�3U�S�XM�*lK�u!Q��$"�*"���-*2+���XG�)ύ+����lQ����{7�Fg�@��r�h���to3����TǰП���{\^L��Y�8=�	�1*���#߶�uEa��[���h�iUy�3���%GՅϬݏ~��W�5� ^��1���U�u�BB���a�s��'w�c~�{D3E)
�T�� �%o��(q���:�H�H�P���a�>�k��l"��旜1ճ_��\��:V�X���q@B���iah� ;�V�v�>8�N�:9�{r�������錊K(�o�v�O�4q*S{F�.��F�H��p����y=����%�����"���F��SR��H�k# �Wno�`�iI�+�p��&���N�3(H�6�82�#B�p��q�UDDp�(�t��By���G��+��B"C���\q��X�0����{�@��s�\������\����I���oe�@u�X������'3�é˛��/Ub���iтzPv4�'`H^���޾KnR����S,�d+2(4Dw+��s(3Q�v�f�+�k�VWՔ �y�?X">��1��=�˺��ن�Z�+�<g)�j�}L�jz����]K�x���6�J0iғ��,��X.Yf?���72�A������ъ�E��SF��	���gW&��-�WDR&�rK(���I��,���>3BްQ��#0���Z��1�Z�2��ٯ$�sT�	��p!�gE�%��r>� �>˵��i$��cU�|	�3z��d��H�%�'q����l4)IO�4��4�F�&x��h��E=�c��k���1F��Z#ŝ鎉��VE�$G�������+.�b' �1�(^]H�&�jB\#%?�vB���4iɵy���}�?S�1[I}�%��t�G�S�V������GΏ2r��d��%B��ռ��ǓhZO����lK�N��=B��U!��1�S�P4����K%�\α�S|bǂ�C\x3�P��*�D�$�>xd��GhE��剑�_��}Cx
�Ԙ8�J�.�$; d+�jgǁ#���8��D�P��\�I5ڧ"�S����}���l��9 $|�}j����E&�qilX���-���T�9�-�chA^r�:*w[�g/����䔓�@y�eNi��G1|#X퓁G�gb/)�~�=(W<��R��qP�w?��V�:�Ol���W�����go�0>0+Q΃:��)�������-�{����˖nJ���rW� �����5�"������s�ϰ>�|���fU&[Ļe�6����,H䮺�d�_a��ML?~GU	��q�����6�#rڙd�&e_+�ft�r"���y���`�Pp�>���$tDiK��׎CUƒ}ޑEn~�!?�;����	�dӒ�O�Q�x�nS�|dB��{Q�������3�������@C�1���QU�D��Uyv6M�(Yľdp�9������XW�p�o��T;���u�s8#��#)���$� ��������)˥qK�cX��зƢ�x�.��yJi.�= b,I?i��u�֜m��0/� ]��e�Ib������<���6�PT`�ʷ�`v�8����7}!��(��sS��*\i�>§C������j�����r��3be?�/�W�'|1���4�c�����w�K�����h�6��E��h�U#J�t�\��m��r6�ihY�fz9��J�
3�B�����`����>��~���ᝡ�i�7\�����ܿ������ ��h0�� Haf�û��oFmF�: