XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��iO�U1e�?D��ߛ����24Ԑ���2Lj-S�U�p.����$����gΦL��� �>KAW�zAH����:^��3���\��^�mAsMv_B�5�������	�]����4��^��0�T^ٸ��V4�V����v]LlJ��D6m?&����DwZ��V�T�Wl�rD�N �i���j	x� +�¯g�(蓯H��k�L��mX�|��l�`3Kߊ��i��@#�S �=HR7`�~v���q4�T�eg���mb���ZFVZ�ݥ��D&����a%W�-�@h������ae���<�w�݋ ��/�cQ4�@��V�H��D|D�;�]�-=$N��5�T�� ��ts3��ڒf钖�Ā'�z$����+���~���MY��,޿��o�ܸ�@H+ĞH2��� �[Nk�/9e#D?ooGM�����ZZ����=�]�*��a�ipM��Ͳ�C����љ�y�I����Y�����z�9WKw`%|l]����M0�s�HS�F�Vt`ܝ�(����Iyݡ�p�V�N`|l�H��U�Nߴޢ�O�s�[��[�<d!�F���FW���d�W������g�41����s�ƣ�p���*�����\�3'� ��d�t�x����KLXU�C�	yf?K-���p��f�Ƕe~z��;-���%"mY��YU���m)�v�l��,�yZ6��R��Տ�a'��!�iv"� �0�_�h���y�.S*�������4�<�XlxVHYEB    fa00    19500�PI_0��O�OJ�Qv]�T*
����@8O��6���@�y���Q�nUz�����y�,%�I�ޒ�� �wu�Gb�iA���M3�P\����!�n#Wd�iP�]E��,�m��&$�r�ͺ�/&s̹��V�!y2.H]EY2	�=�I�L��$0��An��T<�Ķz'ȐQ)o�ZMr�Kʞ�ۺ���3��L����+�n��Pꠁ�|��<2x�'�YP�!u�'1��R��`	t� H��5I���k�����S��̍��BELQ�=ڷ��8o���1�Z|{����H���x���{�kn@���+N��:f��ŧ*��(�*��WǍ�����hf2��r�U�ڦ��e�h�Z���/�⏜:����tx�&�
���� s���c�R��ڍ����t7���F1�+�S�&�^kI�����hG߽���|�9�O��!���y.(-���;f/���u��rʕ�}'�N�ݧ�i+'��֍,����)��*T.t$�9.�T<d��{�<"����K�w�������k�e��ώ\�Pp>UIԢX\2��31{�Lɖ@tP)�'�8��C�-���I&��h�t�)�Ol�W~�E�1��C�����k�F��j��44u�K�xR/
�E�9�}��Y������_��֖�g���Qځ�4S��qP�Ӄm�J/��.��$��e�C�*s1��P�$2
x#|d�>d�w��j�c
���@V�t���������a^/ sF�ϾeeW�z�зPmԊ�[T���"7�혶j�q�e>k�k3���\׀�����B�7jFt���dw64m���*��3�z��ؓ����C�##��--�q�Y��A������ ��������C���t�t�[�[��fö���m�/������� w})l�2<��F�y�x�']��v�^[�0�>�14�H���$��NQ���}(<q��9��"�������xj�p@��)B�b.!E^|��&�G�v��64X���0��A�����<K��7���r��B{��3�ˁ�3��C�į/������b$
#��Ä_=�N;�Ŕ�����H�GD�1��mF���1$"�.�z���6�� M�o:�����ڰ���|�_���
p.�[��j0���u+��mmV*���a�ݢ;��9"�+/�7�BY���ӧB����M�u!���ۼ����9�C����;��O<6�Fc��p����;��pa�qYX�,���g'����4v���ĜE���F�8�>#�^�U�w:���/T�f)���3_ı`���:R�~������2�� ���(��K?@��ا?@�b�n���l-�T�S&�Ŧy��.{q�@N�9�3���$�_Ȼ�IޠK�D�޺ G�YvƊ�[�)_z�TJTf���;����T~Y9���;���%�W��q������X7���K�ז<ܺ��-8�<� ��
\������˻]j�|o��)����*�vW�(�0�M�&���/7�R� 4M�}�����0���ؓ�.� ��S&��B�M���	�g]38>1�GjO$����?�7��	7B����iA3`�m��H��_�j]O-�����T���R�B-���O���,�4�!U1�F��U��C	;,j���|�2������ K
/%h9���(����PP!p�t��C�5�n�N�b��(A�v�* /���u�
�L�3lg�j�� �{f�o����sB[6����ǥ������h6V�4e�p&��6����nQuy�:��+�B_�^����f�VN�pp1r�%3u�e��D���I�N)�Q��U4ub�Q1Y�}�c�!�c���״��
6j�'��58����w�K`.hSѭ�;|�]����ۧ�5]��N�0G�J��d�:R��b>���b<�|,�}|Y��!ֆovW��gƋ=�-�*)�(�d�%�����z�e7�=HzZ���q4��f���CCF���)����:��598�QT.#߼��aMS�h���Dqa�u\>�� �����5�/\8Q��$c�p܏�"�$Z�@�W)�3�b6Ҿ��A6ʛ%�U��ꡘ�3R��T}��C����VE�8�P}�j28j.�Q� m$���M���J��eKx�B�� ͧR��J�ߔiK
�Z�9��B����z2��E����iT�	* �MH�_�R.���L?5�3���m�>�*�ud~@iE�/�u/��X���&��;u�ߔct�O�x��2xҠͬ�&I�t_�	��,3�՟�P�\fVD4�UϚW�m�y�����K5WJ&�����"�j���N�]��v'�X��!��^}K^*u�L}X�B7��G�2�m�k�6c�'��!\�ʭҦ��Y�6[����0*�I(��t��U���K�O���|��s [��h-�{���.:q�#��������@�d��r����%'칥B��.�}}�:%xwi:5]��]���O�ԟ�쟷�������k`?����!�w��,~Wi���]�YŸ0g��^hJ��/����(��O����RzK�H�+���L�D��c���v�7���Kە
�����;��߲�@�L9��j=��m!�4�m{���}˄�L|ĵ���Q'q�k���m�g ��wޮ�<>����7p4"�:ίS��@��{e��4��;,D?O�w�3���K��̌kXʌ�@pQ%.�)�T{�X\za���:�H-�3]��Վ	�F��UW%��L�#,����PI���	6"`	���_+33�#��tm-���Q�0�ǅ����l���̱�	eE�TM1�yޠ�P�	p�ʛSqJu��~=*`p�<(���~� v��ݎ���.�|���r���!5*D� �yHvQw�_<���UvU'G��e���Zp�O-�QJ�� A��
|zi+�q���D&�f���H��ޜs7�0?��ǯ���:�-�%#�z�ci�b�ey��g������+!�&�<��Zg �訆�<l��$�p�p:��N$�Mw�=Ax!}���0�q���_�G��l�g.�"�8O7 �K�JY�T
S�l�RM�!��5mR?ߟ�>۽3i�\��ϧ�k�u�k05�4Kzw����7'�(�ڎ��C-�|6����X:��M������BQ/#z�RQ�ԁs�YW)'�[g�J>�I;=�M��θ�� �QHAC|�Z�jN'�R|�b�_�{��Rck���r���n٭R_Y}�"l���aV���+4�ץ/'����H�	X��>а�J�1||�h]���wRẩ-jĥ'@KGLF���D��7��hI>_퇮����B84���ˎ#�ɀ>[�A�$"{6ǳR|]����������8�w�C�W���ks��$�?3c��|��9�@��oQ�����gs^�ȡ����]^#�G>�\�3(�f��'�z��"J�ֵ73�&c�^��]�qBN+��C�Qǝ��ns͗"�\7�@E�}<�|�R��da[�_@�Py�I�V�on��s*���r�/V>��V��E��G��J��M�:b�-�$`&>�)+�ܥ�t7[��ŌQ]G� ��"M;IYC���̅r�v7�5��%v��~+�o|Y�uz۹�S�^*3��Ň�X@�F?F�ص�X��'�3�
G [,O��n��'�D�&���؃����
FXu�J$��k'�A���c�#,�NMu�W.xVB�K�ɸ��䂿)�U����j��]]�M{���K��<07� )c��4.��;��:E[���"y��WT{m���P���'쥄�
���In�Ԥ�p�o ��!��C��s�fZ��qI3����WG�0�U/p)�J:ϔ���mc�5y�G�05?ɛ�W�~=�d�.�[̎�`��"y�'��,�*�?L�]�6�\hLGJW8��
w�P�N�W_�mj&m�g�æ3p?̾�}���"�w�}�8nf-�j���(�c]��>Yܐ��I��'b<_:0�3��b��~?b鄓�>��8W�I�䈤UH�w��2�Q�J���;��YF�6�����+�D�8\t�B��nG3��G�]i�r��O/���twS#�MRs���n���b���VF�uImF���f4[���s�w��N��u�ʀn��/��ƞҡK��>�iJ�J"�ab�i�hX�t�Ib���(��)�4�9�&��_�L�,�9 �4��L	3f���WI�'%�h���N�v(���@�L�vOd:�ptgn=���>�5�ZEdψ��$r-a)����ػ�1�l���ui����C��[�
/w��҇MǜT-�mF���?8ߧ���7 1�_�C��[�����J�� �=bkߣ%� �خy�O�d�ȕ(8���H���V䇪�~��Ǘ�/7���А�/C�q{M�0;��:��
�Uц�SS����n��e���P��o7��U�5�6���B�}�jd'j���2��o�1�44��Ѹ�&�T	n��/o�?̶_*�Wvf/ߢ�mR���VQ>���o�IJ�A�վd\�ţ�8����9��r�=�Wr�lP����!���?���`��"�����S�1K����3��,��R��[��Z	���,���2�J���#�EM��ޛ�y�Ѻ�ٮ�'��:��o�>�2_�(8��aM\�h%�ն�����P��#E��'M��-l������b8Ac�}�^�cn�����q:������@ط��;�pb��eI��D�h|�;�VQ��׌ݠG�d���� z��AD����8�lM���y&[�H琊7��3O�5Q���nϗ���z��۵B�`a@�Cn�MH�+p'�C�wq���x�kևf�z�Z�"��,�dEQ�{=��iO���Y�@��7F�ˏ��r�1��I���X���K��[���wW�n���O���,h�[i�_�^�Kb��rK#�iN��H���4��5����uзۣh�Y���Aj���[�n���Ey*�\���7��6B/��w��+h��<M�ګ6$�gnS.�Ӻ;&"p����ܘg�\-Β�%���N�C7*{���^[Z��b�4:���!囯��d<QG;_9����}��5�x��S�����0��Y���M���4䛝ɲf���kA��p�\�l��m��q�����5L���+$O����C�
_k��� k�pw��7G��?���B#�(M�����ہ~ú�fdJ�� V��e�y%FnyH��jg���2�Y����]�y�a\V�|gI��U�Fj��p�u���N1�\rpD�������[
�:&�� �בJ��7u(��Z7Ǐx�#����Ej��E������7����ʚ#�U�܍ɀ]A!��Tp0#��s6�t
�idzV`��682�ȭ�G?�l�(��hR��w��d/�G�a
��/A .uj8Z)�l=���_��I��FD����kMr�ř� A�qټi�(��Y/�:�(�����4���i>�M�Z��ky�*�X^�� "������������yW�Um-p/0�MH��>
<��\rSbQ!�[�l�SF7[%�� 6H�s��w�;j�n5����(u���u��]6�;ި�iՖ�G��p
�O6���������t䭺�W��y�ϊ�ѵޏp���ಒK!�d��*��0�����;4^�Tt����#���cR����������3���^��G�m2��5���=i��Q��P�@������jy]ޚ������.��f����i�!���\z]T%��q�͓퉛	��	o��IL})/fC�#˩� Uu����Ð�'���b����BB�3'�^ܳW���c��������C���W��z�:�?۞݅ז5K[���S�ݛ���~e;�\z���L�D�]���8o��� �-�0�>�n��}b.�� X130xg��$f�B#i8��H�r3Јy���l�i�Jd��<�l���#W�k� )�jD/(��<.?��� �PƋ�}$TK��.�mh�^]��c�[٩ �﹟¾���i����w$�~��\)f����<����	|Tta5����c��B�C���i ��>Ry���&+���#�:��#��0��^��!w�Ki����mR�KU�%%�-�5�*شu�o���Z�M'����G�op����j�4?p+z ѿ���ig&K�@> J��x�,�6"-�q��M+�$�KY!������
��aV
�ݿ/�E'��&�"�:���Į�=���<Դ �w�b/z�v.y��;�\J>K�̶Ϙ@���J0���T�*��@BXlxVHYEB    fa00     700�8#V�`�lȌ8���}LەD���}�M�t�Y)B\�[��#��1��(�z���/�>#�%��O�#�7\��\�ֹ�B� ~�u��#�oc'G�遖�5���F
k���a�T�4b�l|�@�`7�dX1L�Y�;h)=5���S{UK!5���c�&���W�˙�֣�T����4�@ZVuj�"1�򽊦���փ�Y��N7��5ӈ�����s:����Ģ�r�Q�����~#��/�\�@�����F�Q�]�J�q��@7j�}c�..��+)�)�<d<�aAe��^܂g!M�S��-����c�6Q�Ƭ+�S�f�V4�J/f<����Dxd�1!�!K�C5��z� �@�HW&���3�3���P{">�TFIU�T$��c��{4s�PH��x�H@�Ҥ�˭'|p����g���6�	����3C��2�S*yІ����'��o+b��^or����l�6j���Q��Y�g,�^�A��ͽ����$W��&[�\�z��}�#�8r���[��U����ܘ��hzs�~a����s�ք�&�2���!e��:�ѭ��%A��8O�����15���F!{N_qu�$ҽ���|��1�t87��AY�$���Tw�pֺĳ�k�>��J��/�p�<����a�j�m�w��:�{d��a{� ��aJ4|���y��-��*��%�dںц��N^�;�w��)�OX(1�2Ϩ��Q0������� )HI���o���F�w��x��H�H*q@ʌ��ݴ1D�>y������&��f�eZ��/2��K�(�[�ü��$P:��4�:�����=)�i��Gu��g�刧j�j�6��r���O�v��x��� ��i?ڥy� �����{&Y45]�ۿg��w|l���x�Oq��¾��W"���-����d 7�0�{��hF?|6��}j�
�Og;������c�x�C�/��t�)]�g
=�>>�����\�K��Kv�߃6q K�\hs�O�ɀ/f��%R��m����n�ڨ�`.Q�q��4}�	�{�mL����ޮ.�]P�GB]��u���a��U�љEy�>�N(8�x�}�}B��լ��xu��/|�aj�_Pt_��˹s�R3N��g��2 �	bh��!�����+'l/rq�g�]b����KKU qM�����ڥ%>n���v��3�f�!Xdbv�ߌ�z?�_^P��� ��~E�b!t��	�rt����nb��m���Ml@�<|� X����X����/*��V���?
��g`Sc����d[+?nLμ��T�1-`q��#��8G�%������6�( d�2��mO��(�"�.�T���U���V�P֞�s3�Y� ���]��×	#dYOߨk��*��ʁ���{��U����y|�����9�=b��'7j�y���D��V�Wp�74,3BޘS��*Mk�j*g/�Rg����XKE��_g4>��n$=�^�3�`,�������t����IO0	���?�CH�8(7��� ـc%g�zsn)Iw���D�24d'�iy[K���|!c�PV�5HB�5��ŕ�6N;TC����I����-	0a��cbjʄ~�A�sHz�x�3�ϴӜCH3uS��(���yz>T�7䓮n<���Ҿ��O��Z&�s�Ty�aqpq����n@͍V�}�!R%S�"YJ?�窩��ޫ
!A���Oj�LvL����i��'����:�$��@x ��{?�Y���XlxVHYEB    77da     a60�[z�D ���N��|���_����Ϋ���d.��*�S��c�����f��\w��,�w�n��F0)�\�Mj=����&tQR0�Z���r�h��_O��[� Y,e_5_�9r�_|=���QE�h��4�!w� �Z�ߘٸK�����L�I-y91��x��Y�]��N��OEV����/ȭ��r��'�-�jE+?)�$����GT�a ��qep�m͌�۲�eT�`�A5p#���������
2�E���cG�~ɶ/<��?ɑ��s�p��jz���o��%!�b=�_X�yb�we��P9�&<�	�	ʞj���Z5�]�!�"��$��=벪:m ��xβ����u�Aj�<��v�M���8@�I	ǻ%d0u��o!��9;����5os-�o8L��=hЄЏ:Z���a�|�H���t�Or�!Է@������y`�M�"�
���M��Jz����/�'7~��p�f�'��L酷�$���@C�����n#H���o�s�t]�oWA5�t�ǂ�t�xft���jÅq8盝=���s:�F��+���"_N��р��%4Uf�K+㮲��]o�1��*&/[?��Y j�;��@[�"����U�Pr�/�����R̯����n�v�(5%���o�����u�����q���WLW1�%`���&;Wd��U�P��Ba�t���r�+�f�CM0�+މ^�5�^��!8c'����|��n1�@�[�metj���q��srO�6�;�5���p��*�ێGƙ�ɟ�!U��y��f�;��f3Z>RDn�& X'h� ��lt�����WH�TL�C�41� ��t&d��S]�k�B89�u�_4Q����JV��������E��yLm��}� 1��)0�>-�>����8�+���������Ĭ!f�'�^�d)�qG
a�֘��+P=���!i�ɶ.w�o*���oKJ_;$QٛŶC�?�K�vKn��u����O
�Ӽ����V%��a݅���E��JU�,�o��u���� ~|;��w�E)����ҏ��l;}��ȷ�l�
�_�(04Ӱ[�	�ױe�e�	�5
���h��<�fڞMP
w�ߚYl^BJm/:�d��0w��M��^;�����8I!2����TZ�phPω����Y��<X&��]M���9_[���o�+i_�D8�J��[�a�DW$�X<J=�|BtW�.�Tt+L�)�D@�"Y#x�,R�íl���������F��x$���io�˝�4e��P�#��R�q�z�wҋ��x�wr�5�Qa��]��ZP��  �L�Q�L�1��q�_ߖw�RU�ڳR��u�r��	�e_�]�g3�e:q� ���(ۆXp>��Ծq���~�����U�/Dh��S�IB�OP���l!I���4@S���0��=X�X�)���i�KlN�S쁱�{��O��T�Ö�,�ϓC��AA��P@�X��lIa�F����CA��Ĥ?���|��w�)��w�ub�fEP�� ^M)����l����'��CY `.Gߺ�w�vo��՝ +�!1� +?��"p:�	|Ǟ��~�K�rh�X��F00��Y	�)��|A!y�l�T�%ڜ2kp5(�-��4{N,�O�FE�8�,���XF)vk*��Y�[ṯ��7��n�e?{��Q��`.�jw��~4�£c7�f�-*��LB�:%�9��)+KՠX��ZbI��/�Bxq>)��r��������.��:��FI�<n�nH�G�ƐQ˂�XD�_�H��
lA�"B�QJ���-L��ݕq3ϴR��w���B�5�!Fl��6�Q6W�;�2�S������Y�qتA�8�����i�H�/{���Uk^6���g+��űF�g�����$Ķz^­X��r�6�I�]�³E�8գ�*�f��9�D�PPJ潺(�G�}-[�gmBNbJ����� �r�:y��M�P��}��,���2�U��굀�,�t���5r� P��\>���Mv�L������"��W�H��g���`���h�M��D��	�`_�q{#x<�`����VFNE�eoA%3zKzq����0)"觫]����²G�+�v:q]`?-vi���<��傀�w�dNyRZ`�O�3����~Ӿ�o�'u�@�lo�	�inE�Y�Q�[}Fl�rr�&�F��2�@�6%���*���ůg=pl�~C����y_7����R��L����/
�>4(�u�\��dQ�4�֓��S���I���#�t�I����4�4W���z��c�i�V�f�>�s$P>�L9������xd롤��/����w%&K?z�����6�O�r�����Ӿ��R�1|�UR��[���X�!�U�1[4���b����X;���W4�f*^���(��������b>�f�C�_���AW�{x뇳,%�ny��/ˣ,�9�f	/	m ��`�J �� ۰w~��(�-05�&��T�9�0�o]�ėB/ʢ��J�s}=��P�!�8ߺa�|�U��n