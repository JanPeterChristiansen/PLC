XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��b�PP��dc<���M��iUQ�)4UMu�mq��E5\^|�^���P�C��B-�1��ŵͫެ� �~T��O��L�Đr��^�K�*Z�u�(ۙ
HN�'��f�h;�f�Mɝ�7Ȝ{7����꿳�e�d(ڀ�v�3���7�h�����Zq۫JBH�rTH~���VKM��Z���L�m!H7Vz����D���#��l���0	��	�����ռ;�㺝��7���C~�9���$G�]:rwA�p� �����7mY��a��́�z��gp��[�Orx�0t����NU2J��Ь/���2��'�7���6��LV���Ĺ��㓲�t��s4�(��!Gx��W
y�z������;^x.���"�Tۀ��,�\��
���I�"�2��}�,���Cu�X[U(;���)GY��5{6Cn�x!ڑ�ƨ��J���*��F����-��|Tp<�,��us�cL0�>
ɫYR6�7���[�[xY2]������B�|�éӥ�GRN÷��P^R�v��o!���H��Q;�W�2�d
m_�x��f�
����H{��lJ��_҆t~�K�V��$' <��1�B�}���{�1)����oQ#��dj��O�#�G�@�H������v,Q�~���c<7�lx�Z��6Hp��6������_�u�܆���&���N犛�θc*�-�x$��~.S~�f#���|��s
)x�_轙�mi���`���qcs�Z2_���%hXlxVHYEB    fa00    28c0:Z������)shy�ك"ݹƝ X��M�����JDRt5���.}"�zg���|��k�`���8�,2?��\p�D��@_
a �i�,E/��N@������L����,�ߓ�\ua ^q�׵|�?�o�7Sw�ɋ�'��s�c��Ā�����ޱ:@_?�pc7��'&�AK@������kA"��~'V-!o�Z�6�5#��(�+��!^R og8	_ Z��q��N�*}����Pԥ��Y��/�{������P����^p}��y���v���_�)�����[�]�#�7#1?��͓r�?Ε!��Ի���W)(y�b�Ti�_��E]����>���H1¯����@F�gfC���,ﯰڿ��@�v������ ,�]�������D�M�w���D�sH㊢��$����(q����f?�Q�#��w���B�"�����%1�N����|�UG��do�~��L��#�Q�:��!�:��E����YO�%��I �5�NmD-�YI�Y��n���t��8���Yd�r��(�
/uy�m�	`�hW��� �ɋ��ɺY���-�*h`^�oXa-{�����&ǖ}s��ʆ���f��� "P8��c�_\�{��k�IG����v��4�%욂�����A 1�a�\�7#W�Jq��C���yp�<7k�����`��3��/�%�'_R�j"���<�,
��!��Rg�~bC���8��q�;�U��u�l*��t�ME���+�p��G��D@-�lT.M�9��q�hOy��la�VV1:�TR~���>��i2fף�*+����JF���R�:��8���	��3�h��E@��ђ�|7!b�ˊ}�z�ٌ�u��5 ��*4����z�F�V���t�z���Tý�S�[�N5)�n�Y2cCٱ�%hk7�A�U�}U��O�qL�~�n�"
TTU�pzW�U��|�o4���ߣ�.9�^��װ�����7�2 B7����%[����L����0��^^�\~zcZ���v6,QCɫ	�"�mD�J��-V�_#��_��p6\����:FK-���v�oE��|� ��#d��}I�m��{A�r$�|�V�E-/G�F��ͮ�u*TD5��*��sO�o䙆�:)w'���D'��[R�]4��������?=!i�"vI&�HW5"k�+V2�{��M�1>�7�嘶��$~�s\�?��� }Q;��\g�+�z�:{
������[D�^��
��ޒ�Z��ИvA�쟡[a+ R�ͨ���Z�I�a�7�4���X���m �;���+3�,mg��J�Ο�u��7�x���;Xn�g����+�� ���P�i�,���8jԒ�ރ$�".Awc=ǅ������D�ʻx]߮�BCK���d�5z��s��!����~�_�����t��r�9����R�g� �8鳯�[c�D�)G^�#^�>LoI���{8��)QB�1�s�ҹ7�v�K���oǨP� W��'�R�8
�aL[�e9�O�/b�m�;��JE����̯�*��^�.��xk�
�ߊ-���*�o�k�9&ӗ^���~�H)J��4%<���\��S�Q ~2��}�0#�ć��2����M���-|���~�}�1�1@{D�Ӽ��!b=��n&���R3.�9Kc��D��YǤ�T(�b����(ަ����CV`{AV�@����|=��DV0�_X�~�Pn�f�$�Nǜ�u0�I�,3���HC�>��_��Qx����-	�Az1��w�������Ц�Z1��+��o$Q
pIw4>�(-��ɀ�~�8w �5�[�6d�(�N�����Z��d����!
�sP(�#�_@*��Wn-Ci���4����M�4��T�dv�-;=�[�q��w�㑳��߅�t����c��>Ou%K��hO/j�5N�a�cXKw���X�$H�����\�g8�/0�S�.�1��%-�+f�������Q`��f"ഘo;��mq��wR/�IP���XB��Og�����94r���T|�C���	fS��3�Y�iב{��Q�b��Y�?Ar�L�� �˧��0vA�d�pX�?\CnX��^ ���!���JV��SsQ��
#�V(f�'��l��@Q.j1|��$�m��=
uv��C�
u+�Y�Ia��?q��@��
�4z(�v�U�61����^����޶3H�U��{{gëW)(ZZ���:�uNN���@"�S����D&]�t��%�0tŃ
��(��oO��_�Y�^#F,���|�Ƃ�B2�R����X�4J`��.�q4��OUpY%,JW�:��bi��yܼ����[���Ku�v�-H�	�����+����q�d�/kik��,���P�G��"�^6��z76D5p֠����p��6Mb�0�ƽ���=��m xSγ�o&i�^o�S���~!r�K���؇Ǝ9�r���7�������>�r^���s?�1�+U.��$������g�9u�h���G�1��5BH �;/_�Ltj��ނxt(��H��<��������ѭ�R/Ə`�.#�@Uq!�R�$�x��h��(��p�P��=���O�����[�<Yd�x�.���'��F����L�"�����V���ko��Vm�q	cZ�&������+�)SGV���6�+*�&_��R'�Z�U��ξ���!)��"+����f�%��AdE��z�a?y��c<ѳ��!L�Ў��.i({J�h���+Y+���U����w]T&�����9�Ӻ����k����-  ��f�"�t"29xoo��.6o���G���)�g�zp��pG:�����~M���;6_~�
�w�� o;����K����ߥ(d��*�$���9Jw-�Xj�ٛ�@��j89���_T^
,-ܩ<����;��?��t�L3��s���:��Hb�:�~�+kb�ON�U��Tp*>�ո�i�Ƒ�f�^�Z��#a�P�}��h�o�,��^/���W#2P��R����]���e��WZ��}��>?�^�v�V��"}�� هX�k���G��8�ӫ�o�E�@j��?r�dÉ�1Yt8�l<UCF���\��N�&辚��I]��h㤉���f���cLM����M��C��G�Lu�k\�`	���S[��5����i�D��?N'`�jʢ�����ڗ�����?��dλ!xtw6b�ƭ��ҏ����u�Pď�b;��	�,�1�f�������s���R{�{d�,����8/V��E�'��ܗ�Ql�>���)luar�S�ʗ�;F&��S�,��I���L�G�JF�\�s,:�A�H���p�����1C�kC���1*�$�~1CF�)�i//���q�$Cn�r����I��w�-��QN�����=�/�5 z�,ޟr*�2C�4p'q�q��u���F���L�����z7�́�Xڃ�&�k�~�up!��nBk�Vt/t�+�+),�-ӊ���X���{S�H��t6;<�Iĵtw��D�\H�2�ۓ���#Фĉ�!�!��<���/0q��r\5�0�3&C* �"���Ot�}�#��g[�.2��)7���ɬ�r5~X�@t�ҙ�1K���.�� ]��Qg�ybZ�@���zE_;����l��x�/�o9U�kl\�8��$K���nP
�7tJ4y���G�V|��wz�&}G��38t���c��#�S����@�#z��jO���D.Nn~���[���\'�QW��"�*fƑ�7�`�Xfm˹�X�5(_�]4����!@x%�^�p��#O�
�Ov�"���st��r�#_n����)j8���������9�Fx����m�&g�+��G���>��)��N�$�=�aC-�9��,��g�.�\��5�t.A&��GG,��(ݚ�������3��>,�.���/�� �蛦�����7eR���KCx�\r�@��׶;y.����۴XI�ٶ�"ʬ��" �3��M���m�.�7`kص�wֽZ�,�@틓Jx�ݿe}�[ly
е�M�.Zg�9#�&4-p؋-IW�֎���i8l�^�M�M��v�/(TT^NZ,�jM��� @=`þ���:7x���:��2�����l��2�L�r��q��}W�6��#~##��Y!~������J�-��Ʈe��ߒ�c�F�l]���{�Mj\_�ý���y�q�4`i^7
=%ͩ�MӨT4�5�ܒ�����#�+�8���S���j����'|�a �*� 	��=q�W�^�@j�Ή� �nׄMgԷ/��joq������,{����bgK/��Tᖂ�ӏT�Y!(�f��XRr�BI�>\G��G����&��A�X3�~$�w��/A}��Y�����$-6X9��%�$�5D)2��]'Z$��4��ύ(���	��~FF�+X��
y��	���1��$��^mA�� �ju��K(�CP��h��;g0f0���&+W7�ˠ�ʒ8�"�h�VD��8Yx�	ۓ�R^!�ш��L�9� 	�4����q�؇�O�+lIo����,�Z�?w~g	s��D����^�f��"������JC�%yp�e8�jJ�'-+��"Ae	�$m�d1��n�� R2�I�/�Hgv�Ը�g���G�4���r^���UUET�	0��;�tJҰ�l�c�H��}�|�ƴE�f�Vs��4^*�����:�GI��E2�����1Ye'h��K-Ƿ� ����tI��"��Y!�`buU����O��5��2h� o�ޟe����Odu���O�-��EO���l�A��> �۟�_�QX��{1�D�M0(!�bx��fWbf�6=_��?<`	�w8W���XRSV_�H(W�dp�U+y�d]w�b�Q<=L)0���*x]	���,��ñ��}�t��h���T��/ޯl����	
�_%`��,���Tq��uX���N�p��'��Gèl�Ĩ	�����	�%�!��oX���T?�A�s3��Ճ�{��HL���#fI�z��A���>��32vQ� v� ��Y����|���H"�#�h��H�ZQ�_h�0���uƌt�'fe~��?�S��6��[�ND�MoZ��*M�i��rdЅ=�b�Z=qA���ɺ�3HLX��I<hЌr͊f�m�J�ƞ'^' 1�RTD��^�L��4؂�tdG�ܼ'ǿTS��/s��bf:�}��=[����A.��LDf�#e2{�&N4G+j'18��jC:��o"�1�Y������+�%s����f�a�m�>qe�eB�4j=tWC�:᜛�@p�
��2��m��v���Uw٪@���Rs?�ink��;N]X�f�e�w�������Ln�a%8�h�\P�h�����cD�g�i�����x+e�4���p�H��K�4&�i�����Rfi��孼U�XU�p�_�f}9����9�*p2�h���B�,�h*�0�	��	qy\$>_b(�/T.��h�X���L�zʹ8�I��cq3���#:JK�@�h|�5$�a�H��i����>�X3=K�(^���5�^j �9�ҵ%�NM&�t&YG�_���dq.[�V_ň�� _���p}������$MY�}�+�П�>3`u�C>y�2dSl��HVx��j�pG7�x����>���vn���[���!���<:�|o����B���T^u�
^�Dc�K"�!mjfb�Z��KY���TS\�ǖ���C��6�N�[��yQ��TPN�g�~E1&x��B~�}��u�<oI��i"���r����Dw[��c;��2��<3�Jg���d�K���~�@������v"���ź�H�鉷�ß>�����zp\�_P��K����Q{�&�k_�9#��r�#�
��зF�&=�G�Z���Q2BzJ��I��ӮU�3�U����]'������я\՝�Ƽ)|�n���;���W�6�".��_0�@�P^o���D��<���ʍ�z�?d�	�aV/����Lz|�r,�V���h��M�&	h��ܖ��hqUU�F׃�
����GџNDJ��Y�Ж��R@@��T��	
)$�g�TAܺVn���E_LQ�W��E�_� Ni�CH�4'01�����LPA%XWH��*���k��~�
:�O�����{���H���7�=*�^�Vu�>��(�q,y�:��+ʟ߶^�̛(Rx \!�)�~������%�N����y����}�ۙ�w9[��Om{!;�a���0.�
9��V����lN��F4 U���?���� %��L�y�:�;�A��T���S�8p0?y�Fm|�O`�{�l�YN�	P΅BE�;��c	��i]'���0��I)�`������d�FC����k����T�Cq^�̯&OX��	+	�r������ d%����b�=���^���c��C=��8�\�.�� ��c!��8�k0PsK$�a�(|XJ�Q�A*���$vMLx��Z÷��΢e��ᚓ�7@�Ȯd^�U�\�C>�lVZf5�x��D��}+��p�L�m��7B�~����CNk�7�
��6O�&ؘ��E&�����>E�X���G�����׺��X�f3$��H�&������O��ۧ/8�;�]n�%�2�IwL���N~���M���c�����w�de5xh�MlΨ5R�.&rc�LB5m/��Uͣ��1c/�^�[��3�&8I@��gA��ߧxg�4�~�<('���9_�6���虖�IU���I���]� �SלU�d).8��[C��i���b^A��z �퍴8�}��4�F#���w0$�����39W��OQ	ܷ �`�y��UJ�:Q�k {����z�9Fي5�|�	ˆ�5��jH�]����w��_�ȸ&���*<�rO+k�G�G@�J
G���8��w���8���w�4HeCowAlk�����َ�f�6j����F�c�B`�������Hh�.��2�8{�V� ��4_SJ S(1)v�墴[DP�ɼg���t�����lש���,���xR��:����y�ܲ��X����V�%zRu�D��m����D��XM��Ӱ���wrͯ���M���δ�E&9u�0�C�_-��ۑ{݁H�/q��V�h���?�TK(������B��y���)��Ymq�n����{��F��N��/i��Ɉ�FR�ۿ����a�N�y ��׍����s8�3��hlQ�F*�W�^����j�	卝� 5����V��L��RXS'֜��+�4K���cGY���J��^�z`�'��8C�$fϊ"����nhK�Wa���[-��1�d�B��P�&��Y�Wj2��0b�����w8:�����9g
�A]��l���]������mI�+������!�Q������#�;�=��i�?ʪN��H��*�Ү�}�$s��y�E�<E�s�
��G�z6�m�[a;_�0O���B�+®ٙ�PpG�l'���cɑ�I����޳��O����Հ�Rh��q�2��E�)�R��%k��,V�+�j˒����
�+,�.�3��!?�P�srƪ||MP����@�Cꋸ�q๯�J.���c&�A���h��sH$a��uM�_A>�*L��v�r������������ɇ��125�"��nE	c90��'�Ç�h��rc���7/�w#xG�j��#�� ��� 
-x_��@,,7�t��޳!1�X�e�h�������N�w'zs�����杪c)�<2!�ꙁHk����T���M�G��rNڟ>r� ˏ�Fz�<C�L���ꯟD;ōd�2���ѹ��S�����Q��1ca2c	m���V��A�T���|��FUaO,=]��٤1v��;ލ~�g�
u0u����W�4�[_�A�q�F�x7�H��	V� �4^�Q�VHU�'��`����;���=� LQ��t��p���p[��3!��̾���-���p��%�֒]���х����-_Q_��L,���Xz��p/���iwP���(e)�P�/!�w����%�~����9��)��l!1Z����v����A�).$��z�Zgs�' �c��>WT���0�=����2Z���64��ĝ@��ux�J����(����T�ܴOLr��+h��Wm��)�9.�,r�y��O�#�(��h����a����e{��5�@���Ѓ������Z�M���*b�zy����o.i	���H���F�bƊ"0���2��6v��x 8��4uyOjm�7ڱ;�,����"����e s���h |��l�Ed7�\�7<���C^f��W��՟� �'[�Vչ1:��}�r7;�=+(t�r�%���t\'�9��ey2�Ό��w��ՂMg��,�a�)��������OV3���Y���s,�ÿ�JV��%�K):Γ
��J&�E��w���dS����9��)0Qz)��x-��&����5�pħ���q��V��<\�{E��v߆0e��3���߹6�`�A�����dG4���'�R���VSK�ʞ��&N�q�.{���L����)M�A�I�8h�ζL6k)���M�v*`7դ�'��7��8���=j����hJ'#�p�곺�]b��c/����D|�$](�!MYT��HX.Hr믉�o��ԜU�Y?����`���fx�wP�K�17:�Р7=�KP�Ƶ�u�.i��ahA~���8��}�U���R�{�N'"�'����.]!zL3�Y�ޱ���'� �}qk��_�*6��C^�:�tu	v���@@��Ir��>�d���E��g�z03?�U(d��7��I)�S��VF���>����]�A���b��F3B�?*
�ي��L��Ӳ�t�WK�W;x��l�G�A[K��䛕�J�OH�D ��R^�]nyRO#�^R��W'�&���[��ȣ˃g�/b_��J��򉒕pa9�Y��TW�n}7*^���s�F�=%VV������/	�9�X�� �(�u�����0�cF���w�W���%��!\9r$�H�0�,=�l&�.�?�T���aB�)�C�b1O�e���J�B!fXH�b�����|W�r��H௧�z�A�@U�1��/S��M뙦�!��㺧?�H͖��WǴr_�ݎ~��:J}l,�`�2�	�Rnw�{�l�+�l��z;��5K���OTF�z��Xh\t�Rkwa;N���AC�� w��n?��]6���7�K�F�ۇ�ݢ�Ç#��Ci��&��M��MBpvRg��C��ܨ*�t���Y�ڴ��ɝeF�K�u���@�y��n}rpt9]��O[R�D�������_
'.Q���&�9�|���p���5#�S�Q(��IM����Q��d
��D`NxiR
�D�S}���A1���:$.%%�pŒ�?��OP�t����I�YTZ���8f�CWEP?3�����5����%tU}��VtA��$�t�\��#
x
헠���H��#�N�İ!�F>L���6�Ww��'�G]o�	=>�>��q�ά����@��~��V~k�.p�ϯD<-n��ed��+F��]T@ߛ� ��7�ig��*��}�Ng��V��R�=G��	� �
��ՕD�J,n�G��$�����n�&����#;���a;v.�� A1e���^���0�@�=A�f��A�k�]y�Q��ɰ��CUR �������������R�[GDx�I���'�48Z��&��u�K��L�S��p�׻U?TP�ܮ�
R����3�]	ǋP`ޢ�2#�d�㍩��_v�RaB�>�P���i5���"-�+	�i�w۟��$�y���K���/�S/7�09T��c#�,0���d���HV
V�i'�e� ��f��ǶjO�:w�����^C��	R�G���M���a�+(Q�����uy<<[ˀ��ϢO��E~�`��|�Ua��؄&Կ�=�xtyTw�a�����p$G���?e_�v�֩h4���%�W�یu[��&ʿ�2���¹2(�g�]���[@�&`�殃��"~�p���؎TϖW>��p�u>J,=�9���Љ��ґ�F�בf��H�S�zzS1|p-��c|�&�B]��A�+��p�����q�u��n�R�D�R_JA��⺩w��XlxVHYEB     896     280g��teÛ��Ha���b4����*6)�W�V>��}eB��S�%B�XE!�y�"�W�K��OU��j]yb��wx:��;����q���X�qXB���t#�Y��,�TߴY(������x^��x��RH2P 9���)���O�bhP8��rBa��n��:<y,A,�"�]I_.6�W��S�2�"P��<����~���X��˦d�/f�3�
��0���gǃ�^�"�����ĺ������i���=~aH�#�\���7��b�ב1H\���+��*��"�,��eܸ<L#�����"q\�1�����]�!m24'U�Md�k(�����^�	/~���k��=s�uqP��~���J7�=o����L��A�y���b�fr�1���0�&���D�&����Ҧ�&3 7�_���d9�݄x1�r�G��&�`��Nh-Yq�H�4�.{gL�E[3g�i�xQ����S�m��YRAds`��Ώ�p�%�%h�O��J��(���O�,�Ss����o�P*<���m��	�n,�_(�l�����R"��If�nw��]��꭯�!�t���������6���w����Y	�co���%Î\0[qt��/�+Ɗ��k�\