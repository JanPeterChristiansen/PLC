XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����}�������BS��RMs��Y�Q�'K�����_R\����<Xї���P�J��_�f�%����kJ�� ��ʀ��l���,"W��G�}�r��x]������L4�=�?���^tah�D�##phoQ��F���P��������c��H�\�{�+$U�����7�(,
u��C��w�B^(*�p8*���)(E��ɿ)]�y�B~2W]��DdD�!�0��F����_y?%�^%�&�eD
��[�K�2�y�8�F�v8;�ƕ��r�K�9$�t�P�[7�/������o�e�BN|z���UL�Ie�̠&��!&tΥ�^�3�d���l�0�Ĵr�ǣ��p��w�)W�@��_I��T8$������ ���*�=�J���KC��G�t�z�;s	�N'Ο��U��{���
�C�D���.��b�4�~%�����i���	���`�Uga�V�jD=���F�
J�8�r�lʈ� &���U�4��ǽIF��y�B����2�>s�=
m�j�K�{e����/-���eh���P�m��;�/i�? l�S�eQHk���U×+0��`E����[���]�Ŕ�Ӗ���Ϻ� r�eOE{����][F�ڃ)�Af�
��Z����p�;��=�O��~�����~U�.^T�M�Z?L���f��(�Y~}�"�t+�kTU�tϚA���eK^�^Ӓ#2�8+$"��C*��u/�bO������+�-�@>�XlxVHYEB    29da     af0�ފ��e����G���&���i�|a�L#kQmqoyL����t+���^ڲIU��'�� �n��{kQ����6�PK�[ ���S�{l_"�ǽsA�?��Ѕ�V�#
x���Nz�&>C� �TI��kw�?�m��{�:Ul[�]��d�HL�-�����]�2S�O���V�3�L���H`}]��ƾ�o3'�y��4�ǘ�U��eR9����6�L�E�%Ca�����;�m�@�M�BI�a�(F��3��i��o���2ZW�Iy�,�1���`�n��/��P����z�ٜ
G"Xsk�c#%�,���]5~��`H��xME/�Ȅ�h��m�b�D�3�ό��8옺?�0�k�R=]��$P�, PFQiTO�ɽ�-�H���;�_��wc�oS���\�P��Tb��8\�o��S�1@���7pb���/|~m�^�F�Kb_���Yu�'x��M+���$��� ��Ӯ��0��4����d�����H�	�Yy\�D�I��Eݡ+=�K)�nW�{zRgL�1u��f�����Rc��<�]�PK��О6�"�!�O|w�6l�[6�Ǽ������^;rtT �cb	~��Q���%�ΠL �-o������w
���f����iŸ��w1epd���tpe���H��pi�1K�B�2�Z�b�)�q����j�*+�v�3�;�4��T6(	r��_ߒ0/iW>�Y��`�B-���qK�6ާ��6���23��(#�i�f�N��V��E�җuẶ�g�|��ilD#��a��POB��v�p����@�J���5W�Vc��j?��tBY����D��b��ڄ���.�c��C�U�=q����[(�5㙷vA?��<sL�L��y�a�-����9�ڠI�1=�Z�A��>�^��K����hz2�����͍�&�a�M�*�L�[z� F/#���f9)ȥ,�u~��W:���  ��EכP4:b�z����z�x�xL}���X���m�sZ�<�۳���X^�^j�V�(�Y�	�.�$�:Ù���T��)���b��1�h~�^��,yC�H4�&|�N�<[��T��rROS�1�!���ȋM���;��+u2N@�׾h4�b��`������/81�Rs����u�;��N�iD)4��:�&��F(E[-�r���t�w���^�W��}E�����c��^;h����JU8��'�D>��$�\z�/����#�$������1϶J�lF�d�^�Cu������E��{��"������G�G�l��q���b��x�,��h}�����M�f��.�ob����Tn��x��i!K/Ɠ(�N�@�9C)�2�i7CC�%f2�n���&����i����|wu^S��@9�:�Y��"�*��od ��X4��Ow� �>?�Gv���yS�WЃۆ7U���?V^�C�����l�� u٣��T�Kh)�A��٧�a�AY�롧 ����{�G?z�f!_9��Z��X���\�c�^��zma��{B��J��$ԛ����G�ߖ�����Ew8���Pg�׃��~��5��Z��^�&p����䡡�1"�T�g�f�2x��]V��e�SO��8�Y﻿���I��7�Q����oh�)�J�:�䜋1�N�Gn�f����-;�5�E���IB��X�ōm
K�#��] L�v��"��f���h�L%���v;�N����W���/���
=^Y����R����"�����]p�I�a;:�a��-���[J7���S���)��)޷11�'��u�ǝ�h�<��ȸn�Q�8&.�ݥ��\��}F}>v
�>D��\s'Fο���C��r��=6��{$Y{�#&�4g{E�*?D���U�S����
sbW�H�T�k��V%9��g)����ފ��� ��6��pc�PMݤ�<z�K%�r��*���b�J��4�vY��`� D��8x�Ƿ	���|��Dɍݧ7윂�Bd�Fyc�1u�3�b'8��W�sJ�-33Pr�U.`�e�g��RE�;��u�r��g�ُ�������B���J���^԰�qߏ

�$(9���$����D(>ey他�3�hk��-���;��*ZJ�����e�\YQMD��*��Y\�;�ۭ�s~7~��*b�s%Q!U���(�����X/[L��̄�$�ik~��C���k"�珶a-�\�K�V�f|K�%ί�u�]���e���PP��[n����lL�7r5��Wkoܝ�yk�����*#n.t�H��rO��-��M�2D�W��!)2�h��������о��h��Q�]���>�u4�~`8��Y�i\h(�J�/��0�r��D�'�l�i�(N�ɗ��":S�4W�Ӄmw���	��q�Y��3��	=B��������%O�(�-yB� ��X�Q�Y�,,L;͵'ҤZw`ܒ˴�5.y@.��d�][Yei��3;I,�JOI�h���w''ƚߣl�f����g Is&%�i��gS��=o�MӒ��CҴ�Z�e�"8�NI�Ģ��C:@5׻������(��H4ẘJ�$��:E@��sSbi6�4��f����Pq��k)�'�N�| ����6:`�ε.�yM��;w����c��Go�Iu��]1��5�[�9F��_ZT��xZ-�`�_6ID||��鿈����j�=6�4���m�e���V��O�6��' IxSe��֓O=�w��.���