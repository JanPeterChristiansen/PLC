XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��`�6Β9��*�}��M�@�J���m����i�\�:f�'����]��2Mi�������"?j���:���= y�X��c&TuR�bܺ:�Y��m��������~g�.ÿ3�� @NL�j7��?k��Aث�ʀ��������ȤMI�t�����<.?W�6�A��@vxN1����I])�˓jy-�I�j�]
3��x�f�WC/b�j�e��ͼ��X��Z��2���Ύj2%�7ԍ�����&����&Z�Z�d���/�^ߞ�o�9� ���\��ފ�0����.�d�w�@�(� �薘���Gk�ve�D>Ԭ�:m����>~ϓ)ɑb��t&�����G�FZ��ԕn�߰��`�� q{�9b9!��:�.4p��)i��S��]"<�.��7�1s���k�W�/ǵ��L4ti�mU0H(-wV�#	QJ���Xn{��yy�5�3�L�����&vƉb���mƤ��b�J���K�nșkb����'�qΕB������k�Z�.��jd��t�h�P�w��fөv��DLli\ݲ)�ءn#���3z~`�7Qǖ�D���;�{Ph�	aV[����g�o��V���̧{�b�����R�r9���~5����ο@�q�S�Wo�x4mg�;����=�,2=C'#En�ueC=�aZBT��H�(�ʜ�D�M��}���r7�en�Z>`��
l���┸RS�h,nF�%�מ#{@:��=��s��CV0bBJ��G��<���XlxVHYEB    9efe    1be0+��Q_���#,c�f��'�D�Q'�YwxC2�Q��*�H�%*lp �лY��3~�PXEN�!�fI�Y���	�z��a1�����=9.x��X����J����H����g��ɇz��Gs.�Y��ۃ������j�l,m9�1�c�h�ƽ���4�ݷ�ܴ�	����O%'��+|����^�$LA�:��k��v���a��q���U��Vr'S��x�
�|>-k�����g�,,�
�QE!�IQ��$RH�/��@�y��&X�'V/�����xCTm��ͥu\��n{P��vk����N8���u^װ4	@ܑ���x/��������I��S5���LF0��>5�h��+�X���\���-�3%��/*2PH�WH��CM$>pj�N�	�;];�1���7і�J�N���	�L�j?��J��J��؅���o�x;�t �t
�5jn���!���_(�߄��ײ��Q��X�f��&�Ŭ��/�8��/f,��@9w��P�$NlΏ�$KҤ6Dq�^�D�ܛ��g��PP�3(w�}����_���Cqa�H�ZZ��N*EJ�y�:��)`,��
u���̈́���}�u�EE��%�uH��_�}�Z.8e\w<������N�P9�0Ģ��-^x{j�>"��*�'B���S��dU*6#�S���%��)��i�NZ��CȨ'YI��*�6xP� ���8��׉���J� ��_�%]G
Y��J$��$��W��gѷ3y�.�\W5���5�[;"M�w�N2��=�F���ӷ��s?��U���O|ƽ���m�n��D���K@g�t���!������1��ji"�'�HIfp6@CUø>��_�Η����e�C�V8�����9L��uD��������T�v����S.+@"�Ԫ�y֒M[:��M����Z��	g��g{���A�f�!M]�?�ۼ�IBY���2Tǿ���J=Y� 
�c���U��xa�p&��b���8 %��v��	x��A*�8y�Q\h�JbZ"M��a�."��yHO�ovL84M�����v��/�|��c|�4�~ >�q��w��L$e5��R��K\�Ӂe5� �"��X�i�����ô���N/q�}D��B�ݍW�)jp��s8}������Y�{Z��t*��v�8M��=�,�.|��b!�=DA ���%j���*���<M2���j.��)����C8�"R�y��D�I>B��]p�2a���A�����).���^��O����e����0�1�+�;�lz����ҵ�n��F\IvJ�4{01�]:&�.A7ȯy�${�����q���3s�w��t��j ~���}S�av�+tx��`*�9�+�!���T����ܓ��=��-F���z+���[�N�X\�t��W�?~p�z��Ks�NO��`�1�u)����zd�Yl��)NX0�>�ϝ��~��[/�_C�K=j�,��{
J�U�E�^Qhg1^�x�sCF^h��Vc�ZS��U��{E��Q������KrI�a���|vxW�]&��5R>�F�T��y�ǣ�~���#�6�y�M� ���?]�Wv7�P�#kG&=MG�����J��˶������ xgb��^X5��7�qa]����]�zP�e��7�MN"��Į��v'��\k����엙�V|9��$&SFmؠ*�7W#o��{�Z{d�Z��P<�W���	W�'�C���s*����6YBq�ڵ�P��=��Ŀ����>���C�;cK`�%�l�׽^�_ͧ�hl&�W4���E�:���<y�jV���/�8����]���3/V
�8,���<���p��]){L����� CX�d�+8�����+����7�W� ��f�ܪ6I+8�Kj� jn3����2A �1ݣو'���m��T4����D��y�E���p狫�:�dc�Q�a�`m�3�>�oY���D%�fޡ�B�pFby���X	�_xD�'��3n)�Y7��������X��2�#4C)p�7<ەI}MI�{b�9w���Xd��@c���1\c�J1�ɓ��|<Z��gh�@�Ɛ�L��P؇���v'����ĈN�q�h�i���hC�&�W�M�B��P��<<,F�툆�g�Vk�Q �E9��q|@��\hQ�]c3X��& �pMЄ�>�[۴�oL��y�
k�½�T�r�D����>�q�WX��(n�����'�8�w�����9d�U�zk�k2N�{?�h!�D� fJ`ڏ��&T��H^i>�Cלʈ��#jF��RO�!L�E��x�&��]�9��[P�����9�ˀf�Uq�K<�bVv�l9�� }��/�z��n���ؾ*,�pO���ha�l��?>��-�4"-!���5��dȩ�C[��܋�����e�F��*��m �1=B3�ˏ��c)������Jԍ@7=4�\������r�^QI�n��Ɔ{�e�K���8i���̈>w�Uh�A����V_�q� 2���|C��,r�%znx�NB�pR-��|�خ��2����X��\m� ��ʉ���fV�1����V�����j��i��+�U�
��'�'v[��ZHA` ��J�۱&�Ū)�1M@�ɊO0Q2zE@�O��4��ԑ����� ����6u����M^:���?�c��� ��n�hs�:;)]WTe7z�jH=_o�+��qd���I�H+F�@_n(/��$���Uy������QLe�rI��M>Y�{��vgnԪ�Ř��A�����4���Q���������;)�bpnj=�����^�P��Ͱ�`�\G�7�t�}I
~��?�vDq�J�[9�=Y�Y�U��rk9Is�p�E��FL�
�Cx$1˔2������gY��i����<ڵŰ%|�:�l\$n�Ѥ�V�2��rُj@itp�����b���K�5r��V:>�isf*��@i��t��Cv�[x؎g#��L�-�-G��/����t��f}>��mb�.䐜��E��Կ���!vus�U>���8��|p��β�jG,}�?���'�w������q�r@���G�hyT���g��y/�5Bpo_�[�M�XXD��?#N{w�T����A�K�V�Cx����i�n5M �<�u�)��S���h����/�.[pS�r7�\S�"���pL���9Ǉ�H���n,�q�.�䍏�H�ZWE�eR������c��T��4ޅƂ�	L�KmNz:�z�C%"�K�df�͛8Ȏ�^�U<R����n��9�k�TL�*�`=�(f�s�7��IX���<�� �A$Zs]X�˾65y*X�3Ph3�Y�@��֙俤� ���%P�l�uȄǾ�����v����x��-[� � �Y� ڣd J7�x �=8�oX�put/v;lp{�K�@�+�dFZt��j��O^�a�
~�<iz951Lx��֧��~s@*���cq)���#�EgA�[efF�βQ��0xWf�(�f�� �I�P���PH�5B�l�7Soɑz>�~��q��}e�[&?ۥ�U��8��ƕ��j<'�ϳ�_X�%�=��qHZ�:��z��)��f��F����xt�x�R�f�̧��k�l�猵��i�c���R�S�87�6�g�p@�id��_�c�q: '�(������"��R���d�i�6��:��]oq�分�^9ԃq[$)I	���\6/��D�'3ږW�ܓ%@/@m��(z�D�-<Qa�k�ʪ�� T9�/��ù.�+S�?xĤt�.wIFc���$�m5<y�\T0ޣW�r�ZB�3��e��_��Wz�$.L��u��y����:����#��瑙x!S���9�)H�	�#4biAB�p]��5�+�8���R����{L�_��L{o~9�F��a�� �9�'�X�g����y,�@h�!�WTG���t�,j#�?���f�������UnUFͻ�{��	\�~L�_1��6d�O��M\muC�)��Ruc{��Y����/[+�5���J�J�P���þBa~���GMz�#�ҧt����x�1�N��H�o��E�
�flN�J�L��o����smCFCjN	0�v�+�#�+.��k��K㯊j�bz_g)i�?C%���7����ޟ�BA�o�Ϟj��Y�" B��o����P�/���»��١���]�Z��y�]v��:�6�I!CDo�2�b�Ԉ�,���fL��&�NR��ş�-KF���&NԎ)�7��yv��o��GЛA�_Xo�fgWA�S���#�Нo��C�2H�]8���|�n��
�C�8�J��N�W�]����{�/G!v��P��jt���zK���D[ѳ��߭�T��f���[M�d�т 	��v`�swuA��+c��<oR?�^f]׍�=�G��i]�S��\�N�^���{7/�M�=2���`g.�&�}6���=W�H����:����������;�NS(��R��wQI���T��9ճ�O��!���.��"ȏe�K3ž
�0B�
�>\�ό����Λ0���㎉�X��8��A���[��癖:��ܝ�����qR�=���f�1*�Q��(-ǅ�mt^7{[u�	3�QMf1(߃(���Z"ܲ�=�&�T{��_��ީy�,V';�h���مT����E0�7���Z	�i���L�Q�������ϣ�U�Ĺ�TE�@W-�B�C�G�/O7�U�u���������^it����Rё�����{4����{V��4c`�a�%aAtdA/������m�@4�FN�FZG���Śs\o
'� �LNH�.8���]�Rݳ= �L ��:�$��]�N5�뽒�kRs��8�@:uV��+Z��_K7�:�Ѡ<	���L@8�S�ZT��P��eV��Ãyh\����[�%�ݡ��.����"'�r�,7F��3X�~t���� +>�|��mb}�;]T�M:�I|����o{��uZ��5�?`�Xmc4��8ۨZ�\�R�=�L#��1�g6Q�޵P�ϻAl�g���� xHe�>A���RS(H�^V�.7?hFꌡU�\>�w:�H�J�g�":�i���ޗ
'�t����Orm�?N���=�ke��k	W҈p�����C82Y�	�ŕ���eY$D8�v�`��$��,��?D�W��B��E�	�+a����S�j�����ǌ��U=���;�5�rC�n�����E}|���׈�Q�p��j��_`�Ŭr+���w���U�O�Π��Sp�	L��^��(k*�7z�ZM�xM~v-�r��s��p�)��Iұ�R�q�O(�K��EG4~�]�rn@�JE� �U9��=�t$�y�H�]6%r�f�@�)b^�&9h X\�R=����Y1�����ۘ��,�
s�';�2����"����~�D8��{�J�sA�ks�:�=�S�;s��<�߼<����^��Z��߽�*Pr�|"�h�rFnC����]Ha�x�5�;7��a��,[<���~vB|�,I)ɨ�0w7�zCZ*���\?y�og�#��\xQ�,�����錥;7M�w�,k*���!'pGp5}o��'W�-p8nD�ai��F��G`fYJHp�v@���HOQVc9T�X$I5vA�ʾ�	��g���>k�@���(5$�f�na���	��D��%���b�G���@_o�k�c�,�[����B���!�gEw[�x-�SB�3|��9��Q/��4���5��!+ԅgC˦�a��Zg?��m"70�I�z�!7�K[z|Щb�}��z�M5l���4���*�ͭ7Ă:K�ч�	Ia����|!�3��Ƈ���E�����e�8��	^��9w/.�-i�-hz�aw;[K.�����{�� ����;O6C,���U(�%�q"ͫ�y�q?."�&s�� �y�w�x�<<�I8�^Ս��?�D�X4�h�Bv'9����h��a���[��0���3.2a�M�_9wv��YQVp
O�6�"g�P���mh5�<���Ì��cK)�~��p�ԛ-��$�/���r�6տ�Y>�,LdwX���Ji�\G ����� U/�A��!��=���j�����%O���z9U�mM�����,�/�(l~�rV��Z���l�MS��f�-��1�>��{�CjYc4rd����T8�!�^7��<�a����#�/�¥���t��JS��_��o 2��Ĵ#X�*q�/EX�0}��� >�U��]R�p�7�r��N���ZF�L��5�\z�K<^vL�'U���������K���28��*	q(B�����/��K�7�B�U\�%/�l&.+W�3��Y���A�pq]`�˷�+��9�������s���P�1.U!����S7���<˜�8z"`�V�|��u��%�^��E�&����A�˟��� V:�H\����z K�p�X6[*�OZ΂��v7Р�=<l��JG°J�f��!�/C1J�mv]�m�%�(& �1�Aj�~�E��'���g︦=�M��4�5�XL�G6������a�#��Y/���B8�}4��c�CT�1����;끮�9߯��������-�n�o��{:<ǻ��f��o�J���Ř�w*�1����.4K]�O.?ԡ�Eu7�}b8���p��Q[�;�E#�mU�e�k��Z�0���h�8���pGՊ6��H��╩4�G���/" ��M�Dm�������� ��)4�#!��)b�{��9d@���?#�D=Kqg������gn;�����7)ȉ3��Õ;V�:�6�vm_G��r3DGLݸM���v)]��$;KK��F�n���ҥ�!6��Ar�P���m�^x�Ud�=�jM��dڧ��C��CKĈ+p{���6�f\y��TsgP���4�2��z��P��56)/{u����N��J�����p&h#�:�i����u)mC�V#���
�d���*P���b j
ȍ�"�at�i�4��Yҿ�