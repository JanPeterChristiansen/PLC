XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��X�j�����~��
��H��7�E�H��?N��x��Fȅ�:R&g� M<׀�,0�Nw.�������
VZ�m��!��:V{���: ����x0�;^�ߧS��s��)�����9|��,����h }���X�岡4�������*�q��	~
�p\�^uό�A���i}�\;i�^,;س��х�ӨH�>���'+�̃�/�װ�hI�PT�`�_"]���8�ȋ�U�^r��z}I�����!~����G�B�}�[�[F�ӒĦ�1�6��b�
��}� a�6N ��S��~�˭���H�#pj�]�����Ÿ$��r:��w�vM�"2���ZC���3ǵ�n�0H���Y��ڋ����)hX��n�̊<aA<t����WS��tp�4���[I­8��X��/��&�e��r��͓'�@��F�:&\���w��V��c��q����,Y4ǔj�)��Ȣ�R�;�*�3�����j��n�+9��H{x�Tw��=?:�qN`�=9�F��@�)Zf�y�"}}��Wwe� "fWI�?v=_a�D�Ɲّ�t������Jj��R������jݏ-b=b>��x��3��?/4,&՜C�t���G90�3�H����%�UT�����>LL`�PG�ӡ>��L���mƿ��k�7j�e\�]E����^C�q3�ph���Vy��щjR@V�WL8�K���g~60
�Y���VH��q�� �â�XlxVHYEB    b8a6    1ac0�_rr_A+b�Jj���n�wLi�2/�x�Y��)o��8�$�}��Z�V���͈Z渿��Wi���A]H�V�4c�m`g��y}�4v��R-
�tWG����'�<�7q�S�}�%F�K�q�\�U�8�_��h�4�;x��A�X�T �	��.[Jn��^��\�5/��8�!��M�ݺf �HV����m}?�;E'�U��)+���i�Ay�z٫xg�����٩9�/����z~e�O?��"89,���)X�/B�/M�+"ƦR2����CE<�	���y��,C�zʦJ�]�<��_���9q����ߕE���>^�q�2�W�׼��7�8D���"~y���P+8%y~�ϢME��k���?c�T��p+d6y�43��V61�F�jbj�V�ZŃ��we������*�$nvdƕ��-,�"�"�/It�7�PD��^�0��4C�����i�Ϭ�"����(ԑ�-%�<���� �a(�f�2\��Ji�=]��5��ە���,�H�͖h%�h��X�z8�����rOt�51^������N�ez��

�ϐ��yU*#)xv��c�5�<ȫ�[Ȁ���a�b��t���X��ꡓE�kL"���ގ�oS�%2���[���� �gsRʳ.$�L��Q�:��'��ύWL��#���ݰ��Y���ϫ{˰�Z���x�a.Ϲ��,��oU���o*��[4�E�y�4E��U��QN��]����6�-T�y�w}I-���]_=
�����3k�pA䂻���"k�����!�.��]߯�و����K�^[#��s�H��):Q$�:�z�T�.��c�.'#
!��cg(�����O:��Z���:�^������sE͞�_S�BXPI� �}�Y��e(w-*�{��e`s�|!��Q�514.���wC���CUϗ���Y7]ۿ(��0��+�{��rb ��u=��Ͱ�K�	b�nKw�^;GKP��R��̅Q�AH/�(�'�m�(��ش����C�?�4�bKKj{Ox�v�9������O��jĝ��שR���k1L��#5�&,_+�}��JQ�D�/��D$�vqO�`�]�����)���T}��-6���r���9i�:u>)F���>CQ������!H4���p�;;uQҩ�B{Me���u�xο8G%�%E��L3�(}d>�#��J�,���5��ݸÑ��/�(��/0�@�O	I+j�0��o��,
%A]�z*o�ϕg
Wk���%y`��Ex��b���k}L��A�tl�ȕ��@�G�!�;�0��y{����`�N����j�`S;|�,u�H�-e_��
e��?/���D��@A�X.��Q�#��-��l�Gz�,��l< ��2x��uDՄy��Y6Yߐ���ZkՕV�(م/9�7����`r�C�]��l��M)i��ZG83+9�n�RM7� b8a����C��K��12!g���1�>�a5�ؿ�O��� ��Y	)!�-r&�x`�1Nޯ���`h�0ݩq3{�EՖ�����5���iJq��4�Lh"Y��fFTp���Ш7T���m�A�|���w��t�����\>i���,�<5�m�]��˶0�YW�8��Wu��F�#�����0�)1 E�<�<f �a:h���Qy��v\��$�L�!"C��7�?O�Y��,�4vإ�$��2�L�2���)�'{�G ������� X�B�y���"���i��M
.q���?Ѥ!� �{xb���Sj&ӭe�:���:�2(ZRG��h��y�^�;�Q����Z%;[d;dj�N��z�����`�@'�ڽ�)=R��w���Oh�$D�V8�n�Z��u�R����)��T�1)�%�p�y]�Ќ-;W���,�"����4�9�N�FnQԀ9���rG�%��ҹ���N[���V�Ϣ�:�˸�Z>&�h{�` 8����8�.�I��x�_n�z�ӫ yX����L�=§���D�\RT׫H*.�,�Q��h�-l�&O���=&UP򹡐!>�Q�_v|-�Edp�ڎ��I�L�E��؆w�fN"-Ώ�y�ձ�[�m�Ӱ�f����`?`_��:x��Wl�h��3M�+<㐏V��d<B`��)�6 �d�>�< N�^V���ۢ�d��R�=����EpZ2Z9�͜
�2�5y�x�(.����VP穳�b�y>L��o���]�p(�{�~���� N��g�������G:!�@qOn[?8�p������ձ��H}�'�����5�5�	�:˿��V�8�b3����O�9��ۊKξ�]�q�)�PB�z8�O%�������>���x�w��[��t���1��M��,�C}������³�t7��4��h�����-��q׽�P7�n'����D�e��u��*G��q�o����u�����Z��샵���E�c����Ʒ"�@j��~Bn���ٰ��V>uJ�l��z�f��ƚ�0g c�����L��0gLx�y���DdX��1`=��řě� 60�Bw��H<����V���Ӄ}{4!�g��B�����iڭ��J>R�Q��~�������bjV��2ߖb��{ŔJL�t���^W2\l��8W�y�QN� ��UI\��E��wP`�ԸT�P�G�	�ˌ���8��A��Uz#v�.��kz?{����D#���
�����0��������9
�١��߹C��ۊ8�� ����}�<���� ��J���Ѵ�^@���������g3�D�D���[���8�@Z(�7�
�� !7�0~���G�2�?r�r���\&Ͼ��*�KN���&9���uPn�wvF�~�HR<�1S��7���b���%�BM^�G
Z��ī�^л7sM�۵�aS�h���ȋ�
M��Z�d,K�'��p�©������b2T��.�?�nO	�0\����u�?B�e�8��D}Is�N`�@�2bs�]_?�o�zL�Ccl�fw��,Bh����8�\��&��<@�����D�Ly���r�)Q=�A�"'�o���*���wř���y�>�z_�u+���?@ϑ@���ͯR�]z2�p��n�Oyto��fP�	$a�OS�����V�#J)�\�c�<�X�91C��(^�u��{y�E"���3L��x��(�6�P����0�o}*,��WE[�.M�S�:$S�T��4�b�'��ƻi-�ap����e�8I\qAL �z'�(7���k�=�(�9��8����BBl�ST����g;F?os*�C�����[V���Ӗƀ��r����/O�k������&�ʏ{�ڨ$r#�yA��HK
o;AĄx?U�d�l��[���a�3��?訥S-SG��Z�y,u����J��Q^=W�{�˳���3�aUGIP�sf��H5>��Q�Z1O���2��!�/����`�5�?4ti*� �-z ��)�`�c�,Q�F���Q�P��������� ��$q��jdYQp��\uw�Z��ި��d��>����B�Ab�;|�,�E��ՆOFf�����~;�#����p̀۝�(�\{��J!v�gʎ�Jȶ�<��ߚ��]<���x���*у��
 ����� v��Ř�Ԇ��)��C�Y{fBxQ�K���(0��9u���E���p�&Z�4M%����E��;yI*���ܯ��z#S�b�AD��N���lE<�D8��]��H� vR�^��CQ�\������̡�������� �ظ ɢ�A�h�-����o�E���vsۮ/W#7YMԟ���{�L�7i}�j>`Ew���SH<r.zG�HS������������1�ʅ,��_+09�Շ��
�l(Fsa��*Y+�X98z �
(}F��s�	U?��GN����D�6İ��p>�配��y^�/�����u���n�u���[;Xs��'�������� ⵲�.M�q�3H�����쎡ٕ3��&/oXs���딥L���?�X)_�;_��j�R�Ќ���[�©��Z�0��Ǝ�Z����ctF����V�#�����:N&u���;E��m�q�ϥ�2��������^S�5���YDn��-�W���wg��s�J�^2f��􎡞Ïʈ����Zpڮv]k]U����&x��@��W�$J������wS���QV���l�#�ؒ3cv�'���J��'���3��Ods�h�ߍ^5s0�^���m�`�?�R�S����î��I3�@�?�����.�MI$d�}�č�9���w����Z��$���m��mB�����&�:�R�}<���ĶX�� Uo�Ҥ��Ҹ9H/`�OK��>�b�¾:6q��CZzWqBw^Q��^��/���L1�E��K�d@}|N�I�E�g�����k��f�.o����}����?���8|X��0���y����cH�|�%lP�| `ҷ w������B�*.W*����k��Oh�q��i*��������!g��t~( f����2z`�69"�.�,��_��vר�������6��2�;_�D���G��Vxz�c�����m�s�9���1Lܐ<�v��|�aD����7il��Z/P�j�b������D��@ �
p�x�v}t=r��?��?'ɥA�(2�Ǜ]Lj�~}�A,�5I������£�I�FDv"�����v�{v�+�O��U���9�?�(׼1��Y�/g�f~�5^�XxI�鷢p̊1nW�6�n��7Kl���I6�k���ᬂ�kK�5���x��a����@V#⎽��<$�J��~~`�D�39U��bh��ٓ�B��b���Q1��A�h�`3C�@w.��mZ�LW&�� �}�E�4*�Gz붛���=?lO�;���c��u]ᓊM}]��9����	�ٔ^�f���!�@��_�	�4d]*�j���Z+�O�o��[���m��@1"Hnͷ�n�{�^˅�
L�Q�{�m�i���������"Q�f6�]���$� ����Y�=�x��?LjLFhkz��2�@J�V�XN��0S�o�L|{�e>��b�p3[+�faS�/��U�3�~SܝMţ��,&�a�a� ��t�*�����=��ؾ1�ԋ�MB��WF^*n1S��9_y��U��i���z��<��4m��(�߀|>�����iX���D��2�F��35!VT?��Z܇�I.�kP�BB�P"P���<s�`8���L#ɐi7K>֓���k�X��B�-iv�� �Q�x�܋��e�\ܕ�4�D�J<�2�˰졞 }�m��g�B�Yp��+N�8a�]��#��B�!/] ����NXR9�NR�ۄ�{ʐ�(�^m��&��~zQ\���w��[h~���ST�q��{[%|#�l&/���pթU��_�,n�����I��Rp���<�O�4����Ԉ:T�h����L����ވ��|������n2r��+��<5� � D�6�u'x����L�1S��R����D@�*<rS�a�
?�'�<���)�/A*p��p;	I����DX
 p�?��}Yo�\��R|��#(���8�	Tဲ����u>�3�4�nA& �
[d�I��@淣+�V(�gO��R�+}!.V[�'#�#4|C~�+�������;�����Ln�n`�w���;t״ý2P�NS5)
.�d��%CU�>�	�+�N��*^�_���\R)eS/6^��R�y�w�1���P?8��'�@��d�Z�[�}�S����$��<8��b����]4p"�@�����Oٶ����0�����}��,QhA��N8.��H�~)��'����o	l9A���}���(N�\P�	3;���>�iHA�brrN#�Lu&q(S�+���]���
��V~E��C0�L��9�Et	8�,�Q�3�52�8�b�2��V{I�L�[���V�ؖ)�y�%Z��[0��a���5h���ĨD���f[<��D9�>v\�V���I��č7�������p��񒧡T�S ��OvD�T�6��*�������c�\Cq��:��:����A/�q��i�8I�G����B�j�x�w�Ŋ �E�)��$�3�Ñ�O��D&*��Ę��%�4d���	>����:�s���_ox���)��d�{���v�b/�KLF��ρ;^
�?1���G�-����M߁��d�K��_gm\����Ģ#H	�~��࣫��@7q=DZ��y���u�J�9�KV��6�T[B>K���Ú��j��ڮ[��.mԯ�1�s�.�r�ؾK#�$�̼S*7����B<��j����	2%w�tF58��[�Vm�{��iNgW�S�I�ʪ��K۱��O�4&7���B�b�}����+�^+el#��k��~dA`�f�����Li�(�e-�q<W�Vt�Tt��1��ln��Y�:����4N��s-�Y���V�$p�s2p���s2������؋�Wt��gr(���<#�Cj�5$�Uʐy;�O�)8l�9�%Gk�&�o˙�Ւ��hhq����� �SIϑ�X��F��*i�O���"*�
�;���kIO����{,