XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������E8�YIe2t�4�t]ӑ�-��zO3�^%;��v�W~�����k���S�Z[��=���k2^<�Z�F�����ːꏈx�a,!nwh����9��{��h��(6E��1��@P�$v�/$��h1;�/1��ו`2ɫ�9N������.��s���q E�Cf�3��0�7�WA�ň��C
&$zZڐ��ℤ���Z��f�G�F��AzE  WO���[Q�B�d�(����Ϭ`K[�p/A�*Sl���E�T%Iܡ`��5��m���R���6�����ɂ%zD�h���N��9������0&�fv�62p3�0`Ax�e��<rF�5<v�u_D�ǂ]U<F�n�̏ �0[_�q�]�.�x�f�P����t�����Ӹ�f��֣W�b��O0A��6�
24��0��f���4���i�)|\_�2e��S���Z�rO�ͪm�ȫ�)�k�^��ȓG���QD�H\��!�'���!�.�"���ӭ���n�b�'�Yg�~�7�4�MY���=wF�4Lw�����ѵH�S�� ��-9��b�z��ҿjո�f������V�'sJ0d]\���Ibs>�%�J�誌���)6��8��JJ�b���0|�`g-B��Jp-��s@Ҭ/�����_N $Ā,�7�e���4���V_���M��%�Z�J��2�q���$\�H66,�������'n��c�<Q��2��؜V�͖~�q�C4�~�����&&�XlxVHYEB    fa00    24706D�e���24�|�}��
��I����ء���x����|�^ƞFo�W�oX����['G�Ԯ�q�' �mȣ��)_ƴ�Ѵڢ����+)k��@#�:4��7ہ=�9���&�Q��j�ф�I���ÝQF�
1H�3S�₟mB�Iƶ	zç���e� ���.uR����+av�~�yw�D!I��?<��`�ASل�2�t��#[Gn\RYko�E���>1��ʓ��E �'�ɒ�gb���yk�?�8��s�Qú|��K���4�Q��v*�ǝ�LUH�uaj����;�U���ZI��q��|�8ö��F�Xy�Ǧ������=�Sm��k�����/���s\8�j�P�o��f����h�c�T�2e�T*�`�c	� �rC�}S��w��[�}թdu�/IVw�ԋ!������%,z��ͣ)|y����)��{I�A�IPp�ܛZ5��������Vk���$q���JE���zEV�ڣ�����1�~`uv:����v䯥��Ќq��g�	��Ҏ�\Y�s �V��ڑ��.�����!d�_�p-p��L�ˀ�N��]/͔t�_[���#$:k-}F���p�/���H�C�y�K�⒳���
�3�1���xK-^�i�f=����?ؗ���m�LQq;`�E��p9Ŭ~��jb��!\V��m�5��%<y�M1p�Y$T"4�`AN��97�?Z�� c��ۂ9�g ��H�M�D �oz}#�S� iC]�-�/�1ԑ�kq����I�d�Oȸ�~�mE�����j�t4�X,���W���^�pk�ooB֒k��k��"�����bհ���y��t��E`�%�3j��_�_p>/������Uf�C�e���������K�(k��Un�0�Y�҅���Js�����J���(q���H ;���]����\#L��Q�iV�i]�*eMg�R�s�t\h	�ؗxȡ4�`{e3�=�	��<����5�)�b��=f`6NC�~��%5079G�}��s�������[�ݙe���,p�
��U0Uy��pV�Ut��T��GA��Fy!� �?R��@�;�
S0�L�8夶���gV�X�(Rpړ �=�&?LjD�X(��e:|\���]]l($�6�A� �o�Y�è�eI�Ͱ�M	j������E�[1lu)w�=#�Me1��a�Ɣ�ۛ�	{d+�βgp�  PU���L����!��T�6���[E~�H�a�51c��o7��MMm��?���l�pv�N,2N��gU�:�`7H���z��D�?�Gɫk�&ިR7,�+��N����~�.��gU����qu]�{��
4�gԬ�z�R5o��b��j�c�F�q
��?��e������,f�o.�b]A��_��d{�����հ�V
u�d��5�>V�G�^U��*x���'X�஖.%h`D&߽�/�;��櫰q2�#�a���`{U�]�+7��!햸�]�r?�~ޅ����������[>��θ��:����y�������#��0*�Ryp��˷�5LU���[u�Oo�>�'�,�e�,=���4; M`dU���J��u��I<��T�)I[������`
UX"L�KR1����b�Ө.��q�Kj=��j~ʍB�#gRA(����5Wvb��lv�Գ�,�(W79��y� C�,o�$B�
������o�]p�J�gκ�I#`^ݖH�V�$z��%�4� �r�o�
�Q� #�x<�u�!����>w@ �#�M�O��[�ö���蹏�^~�
����6�^�LO1;�R�;8j��=��J��ۜ�LK���59���H6�F���2DTˏ-n�1�pH���?� �<.���g���u��uz�Q��Z+W��g�L(E�������c�@ 5�����:!����T������xo�%o��x/g1T;������3菞���}w9�3��S��%�U5+���^}3 ���?��]o�K͹�V`O�-�+ǻ<d�>A��h�k�m,�ZEҼ-�A�ɽl����:�:�� dH���T�_!�C�����R��;�_���{,)�,���r�;z@2?{�(�n�("SfvN�P<2��>1S$�{VȮ��5�B���VSw�/G��������qa1J�%�cM@�� �I��E�,��/>y�3�$c"���c,�S��p�z!��[s��E[/���9dYkɞ�u�{$�'To���N+}�m��R��4�	��W���� ��h0���7�Q[�����]�o��0�B�bJ�vZ�mV�E��@NE����n��t��M��b���  ���8(���I�AS��BW���QQ� ����L���Ji}�$�&�hl육� ���1M���?#Ԡ�M���7$J�ޕԝ��Y�CVx�$�o��5'���=&�t����iu�� ]���J�ii��ٝ#�U��Ox�܊<1�R�';B��L2TWa���s ���A�Z�ʂ�����b��AR��p�ɮ1ɢ�c��n��F�Y�.9��{����X(~П�y���揗���#[E�� \O�����O���SR�L�	|99��܄K��?��\I2մL����O���Op6�iin�{���#��X�I�1��V�cj�;9�hc�F�m�έ��k�r���r^�@�c�&Vlmq|Sy��5{�:dlY�ɰRT #W���N7�g}�l�"��%ɏj��R�fd���~����M�IJ�\�0�q�Vn��tvz9	�9ª���e�q�(p@�3���^4���1�Z2�․�Lo��ט�8�U�H�\�g�݁�)v�v�4�Ο�0ۀS�	L��8v'�N��FM����=�'��=���R�ʣ��_}�&2cCˢ�s��X��8�������3X.N��lkt��L ^�,A$F4�L#ʗ��$�����SV�ʱV_�;�N{T1	�w�O�Ҽ%J�c($���j������ŌAD�0��$����;n 9��k�Q���@,uʈ�*��$�6(fi��v~$|�)���T�I?垿��e�0�ϟ����㓒�b�����J��
"��OF~���F���\�{�^A{,����||tyxn�Ƨ�_ҳiÂ��=�xB?�kq�~���lD�h��� \�Zn/�光�'��[��!>N�w \��}���U\8��IӇK���jp?k�Ƚ��~�TM�����H-��+ʲ�6��r~��N�|.%� �劯#<2��X��n�]ᦺ �xPچ*+�_�������p,�oPL7\���8Z���R�8�K8nܫ4LD&������O�k�7��q��y]0@�E[�iu�[6V2��
`���e'�q�YӖ�>X�d4!X���U Z{d�s�`�E17ڊf�4�-)�ɵ���Po�}��҄��~�r������R�Pz�Z��}�aÛ�?�ȣ�v�o�%ȒH���?lw=�`,��L?�)c��YIi��0��p��O-�N=	Kg��iQ�[���Y�O�F��i3CEv����\������z�v�e���F���轛�����X�~�'pX@�s�ld�z�&��a��/]�����N���/����Ý��;k9Y!�� {ڽ��Ur��I�<���{O��A�
��� ��E8뎳Ի�_^�^���4x�.f)Ų�������������������@�&��V�u�6�Vُ�<�lY��Z<
L�3��[�Ǒ� L�Pq}+УW������I��^�`���'U�$�y�$�Q�H�L��1���k1]f�MѠc����2hd8�J�,#K���L0Բ�cZ��"j�JB���ᥰ𺉸[x�v��w*Qǘ��u-3�M�	�#i��ɾ<IE>������m��zɊj��N�y	Z55�in�iƵZϜ\�E����X�4*,��Y�8PH�ꅯ^�,�x��S]o����!���T�!�;����Po����EG��q�O浈^9���!�_a�4e�	���%1��մ�W�CہJ���q�$�]@jA�\�~��.f�+�����~[��y��6R�%�� cxOB]u7~�L��B��4]�[>iwW��Ԍ��<\0w���k�҇eQ�Jx/�mhY�G�;Y��� �����);��
���b=;ڬ��V���o�T	�ރO�线�!��+�z8Xڼ��8g;r�@�׎E`���$Yf���wsG�h̩�=md\�c�"@�6}T�e�!�S:W��a�{!ZӠNޖ�C
�{rۄNH>���~�T�J�g|�r�iw]�p�`�g����.��\��]B�+�}��y	��)-2Ϳ8M�uu���Y#���D��p�7���]Y�� #n�rc�-"P�FAó�1g)���������{�����g�B�#KPX2��s��1����(\��w�F��sb�U*$��7U�m��fr�@�y�bb�"-��������\�5T�e���qa(�ǏK^�f�z����X���V-H��0�i1=z\�[�{*,�A���0g���}#&泶o�J~����1Qr�]��i}@�Ҙ���Z��!�/{�'G���O�p�?��з�y@A[�3MX9������d���ie����HY0�1�����Fw���|�9M��`�e%ł"����y�4�(^>�ߐ{. ����P|2�.�r�o'ۇ�&�a7�	�fo�Ua}���#:ߎ\�Ju�H�Nv��@Ab����
�yTK���5d���a�9������'W���/���*WNv�md���`��ƘF���ѕ����ShM���|�%d[�@�`�ad�F[��]RcWe)�j 
�r�{j�|�h��@��Q��Y~�ZI�*�`�DʰRZ�$� ��g��/���{�~�q�4W�OI����i�g��b�L�n��A�I�� ��g��Pw�<�PZ�~��~e�%���p��R�s[�}x��(��ㅥD8�UQ�V)�N4�����������y"���t�C��,�+�ɰ�Z�5xx(���� t�*�ʢ���{����@���)���/�#ꀛ�5��cl2���p���#|��y;�W�	@��8O��$�hk̘��\=wskl(u$�5 �ݑ�|�����;A���ZZ�����	���~���4��.EK�����/ZO�1gA�64c�X�3FhN'�+w&=X�b�Y#VF�<����dk��v�^�𘉛�NKÍ����/��\j��ٸٯ���iS,�?9�E�w��j�Fl�A�I��Q�St�����4L���G���uǄ���G�.�A�·�3>/�I����`	���f��������8b��h[��Z�bY��PD'��e=�����pG-��ib.��3n�j�,�Q�=v6#NSyT���
�jH�kP.C�W�ӵf/_#���>�Y2���G�N(��+V�n(gR��$ ��_���U�X��a�)d�"SS"\���5@La����9J�H� ������x��>~������m�>�g����ʁU�~����E;V��3���5�d�+:��T �8s��v�6l�9i�y����N�Eꤊ�4�kDN�v�&!)����	�s�Hm/J=����>�H�f~��$%�9|N���a�Q���s�%|�@�ypt_G��R�~�0���"�۶�S �����Rx֊�S���C&�a��ɻ��	��*�ǅ��G^��5@@��1�%��=�����_���۪FI���%��_���.7�X��3cǂabK������Z�ʭ)h�����q��O��Q�f{�܏���@SX��ݤ��
��y����ۦ�*`<ݟ��N�.�{*&:�.�B����t"j�Gq4���KL�)N����M���-�У��`�Lqȥ�+:�\0^��q�D�A��&��Y�s��{X�e�����P�ۼ��nnG�(�����Ø�� �a1�#��`�]���4 )����M�4�ǐ%% �B��P�^��Q��N��(yA����弄����cu��/쭣���������iH\
q4�6\_�z��x��'x����0mA��#�!���WI�w�@�q�#L-k���2��4XTIj_�y�K�����,@��< �5�OL�%}@Q�`�p5ϝ��Ծſ���@Mf]��&}w����4����MXQ�d�C=��� ����>���+���xAQ�آ�m�V�u��W��LNe*�Xpu��JO�[5Y~�S�	J���5/ej�8Q"��U(�ϓ��(��Ƨ�|<ݗ't&t�,�1�~ˎ�|+Rв��S�%>6�����<b��m}����;������!�HWuoa��tѽu���:P���ВJ#1s4�LI,� ��Μ��`n��m��@Y��O��Uz����I:�!�?u��	��s�X�-�.ηm���ҒtD��!�G�3u�u��9=e�����*�^)�ԗ���xA9�N[\�2��jK����?�t/tD �	W�ue+Z@�$BK���H�	�k�DW�t�V]���{xG�]x��n6���̜ 1Z��Z.�Ȅ���0�2�tS8�`�/RE����v�:
�)�������[me�6���PfJ0������H1s�?�ev;�Z�$�vC\�����ic��:�|�Nz^(�;	��^�r,��F����Xvǌ�ɗ[e���V��X�����(<��`LP?��w�=N&��>��B&�7��W�u��9��Iw�_�.�k3�m@�	�%�%�[��`;Q����Ir(@�c�~�#��=�Lԃ�$��G��$���J^8��u�UUp�R\"��d=��Na����=N	ďV�l}/=u	���z�n�(UT"?HL%0q�,�A83V"s�E��Ɣ�*a�j�:���=+�n����a	6;%yv
r7��,��QE`��d?�Z�]���J�/�K��wM��a߼�ĞBa����������)F=�$:��KK�Dا*����$��[��vS��E�~3�v|��
"����U��i�_�Os�Z%X�� K���:��nr�]|F���4��˯ʀ�|6=9�Ƥ�x�E���;uyHf�.�TA0=�gri�pҸ�%=��Lv�F�O��3+�cݢ{��dԾRGu�Ύ��-�yUu!L�b� kVX�����`b�f��_5��W2.$�������T,9!K��Di��Q+?�����F���25}K����ۃLv^�.���Z�>$=��?��ӷ����A��� ��Ī��bH���p):kP]�5RҲD�\}覨-Kc�]Fߩ�.C+h!^��>��rs�w	�~�@'o�+�t����;�<�l\� �WU�Dj���v��)"<KƵWJ�b#[�4G������-xS�*��z��)�����J}��&>6&� ����%ߏ�p������iU�\V(��$��͊~�q�[j��L�P�9Î�۹��'ڔ�-�.���K�[t!�4�-RA�%����<N$�Đh����GQ��o�`��G���*\�k+�!���X�;U�̋��pPN��C��X���{Eo�٭�k�"�_��\�9�G������j+�d�[�%	��MsS��e3���
lS��6�Yh����z���3t�$���&V�p.Y���Z�z��j�@�G�ҭy�p���x��60��!���Q4XS���We�i����#��_�S�Hy�7�A��p�K�%�Uҥ���]��7h~A�m��?�B�5�kǠ���~f�UY�0 w9��u�4���$bJ����xv"�� >��.r1��0~�H��Y�ˋ3�P�L�C<wl��h����؛���<3����A��¬I�@��{�ɏA�%v> S$��D���q~�~�T=����<l�+�d��7�i��3�y��%)��ؚp�퐣�-�:���x�����D�v��,.F��h�t����O�B���/�X}4�r7)(%���)�&NX�s���J�Zl�??M`��\-o��|��|�6C����뭊��������IX EB��5i��#B�pd�Ȫ.Gp�jZ��R�W�~�u,��h�Ԭ9�F�������V�4�R��J��5�\%��O:���Uj{;��uo,E-��&�v�u6�g��L��!�m�J�n�H^�(�]K�����L7�b���W��fah��";$*E�(hb�ñ���jS��84�4Ing�*����
R��y���F�"�٦�!��E<�@�u�qNqm�H��\����$g�:�a(ff���(���eOnD��2ߙ�J%�9��˔[�L��.�#De�4(V\ H�����7S�7M�D!�
�n����x`���|B��#=���<K����R�Z���vl�o,wD���1�~����gaQP�G��領��ģ�5%R��M2yf7�?�Nٯ�������<�Re&��I� LI��&���e^TU4v��_&�,)f>߹�F%��� 0��_B�,$BZ�M�p��*���7h��%O4j��̬����/�G�H�|�g�P#S(	�T�
���g�-Q{+56���!��͝�`�c��.]RO��.�-jM�� ��w�Pi=����G}�y�ǆ�������[jEWy�?+%��{���2����/�ݎ���7�knK�%z70+�6�3��s�@'ԇ���5(*\�nd�GK
�R�a����� �g�ZO��ܚ3C,'�(DG-'4�<ݺ��֤b�43o���m�JW�VD���W��,��Q���6s��X���r��D��y�wV��;��+^7�bG�B)�+r^Ȑ��*�g(�c��ѯ�(Aw�)K�D6�l�c���+�%&WqA�uQXZ8����I?I���# ���훤���K2'�R��� ��v���R�CM3�`����{g�h�m� 5�+h��a����@²á�7��nklJg�D����%���J̋�vk-�{�[�(�D�v����eM�q����%�R��G��d'Z|���`%y(��!LVR�v�_"Z�忒+�\��U����|�E��FE��xcK1�t9��3C7ٛ��8�c��kYQ���s^@�˒P�)��6q��.�.8;8��Vi���w��!߲\�گߦ��/����%^e����
��S�XlxVHYEB    fa00    1b30�IAx��Y+uѯ���̜���穵rӢ�s��P����Sw�V��Yr���]N�K�Z��S�������5K�WKF�d��^��,~�ӎO�5��=���D����EB.�����vm|j&��c3pw���3c>��`[c���}Kז'<oA�(LA�8m�\mT����7�.ڃ��"f�D��oE�֒�a�����˟� �/!(����%�m���Kpǘ����z�l*V2�J�N�cb:��d;F���0#~�RD���j�6ZzT����?�9��v��J*�u�J������>\G�l�r����_�Fw	RvpW@_����`�a>&������ixT�]�� qT�E�0��g2�3�  Y�4���o�ǋ�Ð�u5S�A5������hK3f0�R[�G"����V�p:�l*��%ǧ+"��rI�	΀f�/"�"OZJ~7^�߭�L��w(d���
�i��Q[��[T�^�j�"x��M��/�cߵ�,0bH�P+��?�P�-�`�|Qҗ2�y�Z�b.Ny���\����Wƈ��[�!�;˧���I�������t��,_�n8 p#���\�x�L9�:�I��ՂS��5AV{�/>���ec##\]b	F���ԥ�}�kN��q��+�5a��Km�*��~݀C�6�>LǼ�$Cӆe�^�(�G�qTz�M�	��eD	�8�ީ���V�wY._c]���7�e�E}�߇&�󆔴�[���[� ���㛝��)u����׻���($��I|ۆ�*;�p��Ӵ�����j.��p�L�A������	�X��RB�W���(*�jƑ!�gt��-��E�xE=H�-�($A���Ϥ�b�nMOR�����>��5�Mͷ�X����[b!��@u,*�_���p�(`�L��q���(F� ��9��t�R ]	���"2�Β?�H��+[���a\���i8��7��_&��Q�3���[u�q+n@��Ә/z��9h�.	/oN?
�S�q4�"��5�w���ze³���M+Hu<A��|���p%Q�����'�oG�L���ȅǼ-��Ʒ3�>�д��D�E{�>�4,�8;̩(�R$هw(~
���i-��2��?h�[�7�2+��3$��/H�(��
?�7#�tB2�n}h���s�A�G+ ��Za�N�I-S����ag��{;��'��fZF��%�&���}��_[(k�scUi<ݰ����5�(���Y 1�3�������� �Ƀ��	 k���sk`P��GK�,�[pʚt*a�c"���ѻn�QLȁ�<�E�PV������%���ԣ[�*5湲��" �_.�V�/���D��[Naz����6����G���H��VԱ�'�G���0�����y��=?�h�kPD���8��&�9\����s�A.��ӧ<��:c�
��|UPZ����NK3���{tI٩�@�}��B�����w��.2א�k�UE.���v�}��d���O��U����d�2a>�$(H��n���9˧a���Tq�����+f�&$ ��8d�C�r��T���u�� ���҅�13����$ls	��.�ǧ1�^���#��g��M�ߎJ���Y�:��M�ل�i�`��!���+��Uꟊ�|�~`�	�`l�R��)��Z��Zt��ݥl3�\�8p*=)Ld���.���ZH�4yo�"j�L���5�d,� �a�T���W�U��0	�&�!9�qUI3��o}4b5�ʽg�],8qC� ������=����u±�ޗ�ey[�` ����x$?P��Y/|l|�:_^�
��8�c�� B����x��1n�����c�;�Ԣd�z��{��9^\�潉�@�v��+OI���5���x�7�aj;���ʗu�{K0 �i���$>�h��y��u;Nz���j�#Q�PCe�/!`��D����nFY�ߊR�U�8���Nq|�f�Fć���Π*tK�'i�n�!����v���s˂�4#����������m�s�1Se�ܒ�$]p=2�]��ק���tPm��2�8χ���"��S�Z���Kz���}�+|R�C��� /�z����e5��Z�r����w(�y� ��[�ns�Ѯ��������#Gp��u��B?v|Y�h��Y�}��QX�Z/���Z�;���H�Zpuy!��`>{�La�Wv�l[�]�%�eOє�b)�n�)�CegEi�B
�1���/�k<�L�7M��|t��r~I	q}���=71�☀��p�.�����a����$�F3L�*׮�ca��\eRűd��^]<�;"�y(��T�)���ș{\_�:&S*@�ڕ��9V��_�h2;S�tb���؉�8%������AV1(�[����
�{xK�!��J���)1�.���5�U8a˔�g�α9W���
5ω5����u.�T�V�)R�5O]k3f���؛��?}(�2K�-�w�2aF�:-v�\�ؽ����&7�N��o�h}�Tՠsl�[�nfLL㞜�I�'1Ӹ�S�#�鶆*`e��V�z�ֈ��kI�/^7п'�8�`[b%yٿ�Y3ZFT� �t��z~��gM���?0"R���<(�T�/�3�l�:QT9��*Y��Ik_�i�8�c�A�a_(��¿�i#�q�u&Yܣ��ė}�R+J�+l�dó� �b^\�!Cm�Ϩ%ˋ����LJJh}�?^~��ďu�a�.DVb� ��{���|H�[* ��Z(U�j�O]�5���QI��S�g��kA��i���rum�9o�����{�cʗֶ�k�p3� ��·f ��儢��B��:��������F��iO���,���<�0:���!;>��IP�kw1�X7��|J�j��`�} u�K%nN�w^);H�l�u��w;[61! ��E�.(�4�M�'&���̏UyF[�x�4�)]J"r�יMT9˼HÒ_��$�<U�_��v�s��5���J�����f�'��Sg<?J~���~�|c��-���LU��Z�������-��_o�U��X�����upC �b�:U*�t�����}z�)�^�X�x�Ӛ)B{gn#U����]�D|���+���T3~��6йU����_�~��������K����Zue�L��m�ڕ���z�cI��`V�Z��m�H�b�n��N��.�>B��B��}[���+������(bs�s']���]BFo��hiKԗ�lA�
����UÂw�d���:�Xy�������TD�8��]C:�/ʯ��h��%�pf�p_��M���t�"�6�S �[�.�]��̖�� 6] �I����Fc�\tN0q�b�m=�����=���x9�"I触�̻�<��zg�+���>�?~� �Ro
�
n'�$�Vn�@k���R�%����,f!.��D�����%V��ܾ/�����o7�����^� RSl7k6���ze�@8!ML�鞅l��*��,���v�����A"L���!W��MG�yZ:f/����v̓�yf�M�;%u�R���X�Lwnb}�H��M=X�����bW�a�9GT�<��}�o,/mCB+��YxǊ�ua�9�M6�7JR!"_�8 o��U0�}�k��0���ba/�k`n��N�T؏�>�v�>��<��c6��*���m���]!U�����/,@k���ĳ<t��=H�R�#`+ӛ3�����Ǐd�cuؾ����Akά�k� ~��H3�T����]R
�Ҝ7���d��b������@��	�$
�I��{���8��R$:� F�[��c��HTV�p�>�ģIK^��]n	�V�a9�ٝ���(ؕ�����M�����݅v��5����LF�9^6�"���-0��.�/X���32]�{Uo�jS�=���y���d�d�d�.�Ց��D�Qv\�<ni���2 |(�.	c��Gx�0��ˀ�4͝d��P��ܝ?5��L*A��t��F���4��C��<3���j�v1X��
��<��(�W��c�⼛�׸6�t!Vʾ<�_,�li�v�s�����PtHwqp�.5��0�^�����M9�P���{��I^��0���ْ�lt�#��{���>PYqS:X`
��x�2[���q9��z�IiN�����Z�X�3?�+�>�c�����/O�NZl���C��ݟ]H�`�1��ڶ7u�����o�S��sR�))���Ә>�%�M�����r�L�F��v�������'f�S���Ϭ<lU?�ЗB�"ŝh_f
1��$�e4&�w��S�"�����w�~"��x�-�������nhg�y�j�7/T��j�	�E�9Obèf�11�:�פ����l|5eu~�\��	WsI���LjBZ�:q񇞽,r�hSB��l����F�`���&���J��ǱÜv2Z�?��P}�Z�"&���/B��*3je�j}yejI(ꑋfL
���%\̳���$�%�Q%N��_�u�{�Z
q��,��ໄZq$jT~���e�>��/|Ie+D�
�6����VC���{h�ƈt�^
�iȨSnmⲻ�{~f�_X�xp�	5������[�Oj���#Ø�)�ϼ�Li���ک�_5Z�����C�KOչ󽖓���ev\s:�{�~��]�26q_�@�[|z6��Bx�ͨG�`�фO�Y��|��.L0s`��dp�-�������z�,F#{�o�$2�"OEC�k�9���U�KD2ҙG���(�f���פ��P(�����;LQ��� !�v8�v��[��/�?ޟ2��ѣ���Y2t�'K�B���<�+�}�-��Oϋ�pە�޴��)Ԯ�oCH	�_�mw�*Ϟ��^Y�A�s��"R�@��W��%��nG��Q����RL%.�
 (����ŗ�''Ψ���ml��ӸXB��c�C"N�x�/X�n�:Q���"[���kU �p��/]r����!$NLfy�>|�NE#�aX���C�/���̌��yD}U�D��\��(h,��u�Xn���7��/��>y���bw9,�&>ۣG| �V�Xk��}� ��_�xU#��'u�C��װ��$���f�2\]�u����"{�y!k�o���Q����a��=��Z��	;|ðK�&�ܣ2Zt��f)3�/:c����D���Ӧ`�������b?�_��p5�\4qqƓ.0�	��I����Y�A�6@���[4?�����NzJs���a��}�C��Nj��ksǵz�\���F�ݛ��?�������o�8AK�#��R�62���<KU�0Oa�Î(ԩ��3�\������g�wTS�T����i\�!�)||c�R��I�(�&Tca2򃽮W)��p����ҾnQ�[O>�"l�4�� �+Y��۳{.O�)��k,4�;G˾���R�5��~������ٙ�<(�k�oq�:����g���e��J	�U������b�.8�Nm�69<"���~
�I|���3�"�|����P�?އפ5	J�W����A��G>�M0�p�0�l"�i�~S,.ь�! �>j��� �¹�I������2��e�o^ ���׆��:��µM/yDH�3��T���~��B�:w��f�V�����=����]�%oi�楨�m���Y�w��(2.!���+BC�"��^Lv (
y�{6�L�/,����X��.�Lp��\���q���q�����Ԑ5�@'�;sU:�׋�Н��ÕX��/��NI���i�z�54�L��z[=�1.���(�k�XN{�e_�%��*�qk>b���W��h�|�s��[9^�ڨZR�.Wfm����j���ro��=n�w���G��#S@1g��	���k�Ih�n<��)�>��K�D�_+�}�������L��fO�!�y�=d]d%��c�� ��Do�C�3��J�n����gB��zR�oH{�F׸��CB*�&}� zcN��K���)���T�������:dcZ�B��P�"el֣SC�gB1+�]^�R�C=1e2o�q[ok���C��`�?�V`���X~>���}�^^*E�#��e�Ӈ�r0��(d9��/V�� x�f3�A 	��,L��~!1���~�Ҏ?3-�s�ϟ���U�f;���lT.0d3����W=��8�	^�sp��POHx0�u<�>�E�]�����Ŝ��{j���!�nKII��7��Y
����&Za�ju��Ip[�f~dߎD�NED�ڴ'1OU��#Ja���ꋌ$�'�"1��[�!l�4x���q̏�)���&��-|}���o�������ۑ�㛅�]�N\�f]^�T�\�X��l+�����o|��eSQ��C����4Fُ]����\�7v�wV�e�7@CV�����%���"��2�,h��О�Ť��;^��,��oR�7O�r�R��~�����Tb��Ց&"�B>�y�����f"V�Oe�4�T�������_�(�A�Sg�`��FT��${u���ewտ���d&m4��x -�ϖ2wʓ0g�������Ȑ����s�[R��vlj�2��*i.���V]��L����%�]2B2!/����Z8"���(��c�}�a���IR.3��טd��������#~&�����Y;C��ڸ����I�C��}X�)�Nx�{��J�Ի�)��|��w��0#�=�೧��1^~�F>��Z�0�����Ƶ�\�k��q���c2e�*�1�%�XlxVHYEB    fa00    1950_V����-,n�v��L��s��rt�A�^lU8I���n�e�0M$�Ø��j��y?8i���(������f3	z����r�p��J�tIH�=�U��}��G�ē��&�Q�#k��[8�P���mP<��G�Zc�F�h��{�!p1:�O�"�z�.�t[���O	��H 3�ƛ3�x8������o�x���kCr�V& ��`����� O�V�Q?MI�VQn��7z�p�x�Z���lhi��Z��|��0�ʨm<�r��D��H=^k(��b���4F��j���@���8��J�~�h!϶�= ����y�2�}��k�?	�퉘��=i���F�O@;�GTJg�񼶰3Ǻ�a�(�z�a�8���5�p-xBj�>v/���L9��e�� �au�}��6���թSe���<#@Z�p�x^F�b�_~���L�o��&W��c����7X�c���D7H�~")a��z�bh��r��W�`*�i")`4H>]�Ur�;�5TY�^��f���D5�����ۿ9�_��O �j"�� 7r'e,j�"H��8�!a�b�W5�a��`?���2�rR��*@1n��P�� {db��ξu�����a^%n�o���/C���}ZY=���ͽ�%�̥A���'�u*+�s�k��������t�&_	���n]�$����곗�f�SR]�m�6�O/k�n9�����03	I5$0,��P��'0 �_�?�E4����ct«|���v�چ��Nl'��z��x�W��@�X+jSś:��q~�WtA�X�qD�&m��R�N�������:���9@�oޘN�ЩK�(T��ڙ�T�ƚ@���2�d*Ԇ!�Ɵ�S��r=�?��4	[8�JџA�{^���;���΂�@J�<A�Ihd�*�
gA�n=����^�eO��������d��ئ.)�v�`ڐ)��)�fضL����K��{L�9�e�c�y��,�Y⨹��4-s���f�:Zx��/�He$�k�V�F�8��X#��d�쬵H�3kr	VYD"H�#U��v�b�i�4�Y�[�J-�B�V��b��	��	U+Qe�W\�fFEY>
*�l;�i,9�#����.���iR7�d2�i��x}�'㥂)6.�hw-�UHW���#�w~��%�V ��f��7B?zth���og�C�T9lK�8�cIyF��P��{����Ub$��
���ȉY������k¹��_4_�-�-��qS�+�ȱI��5�� ��PA�Ȗ9L�N;t`���F�����9f#���w�����*�':j�>�qݳ�ޖ�=1������hۋ�Bl��ڇ�g���\Ƌښ�6q��QI<xڲ����ԭ,ACͺ��/M2�+m��	h��e��{N""ncHѝh&����'졃��4Kx�!*H�SМ�gJ�o��W�sbK�S�T�\+0�ٍf`!-d���2/<Ij�Ssg��y�,+U�c��{G�����7m݆��'��Օ���%�;δfc����>�嵲Qc�Uz�b�3��­�����?��kS���AK�yo�o@�  -U}�����{�?w�",�p��Q��+�۴����C�_�%�
�הLX�׺i�Jt�JqY4"��!�Ѐ6�;'��g/+\���5�Ҍ��l� ���ϙ�Pn�E���Y�=�(����C�M+���E#\,nv��SVv=�Y7m��y@����t^	dI:?��8XNW�{�hs�SLmR>�* �Q��L`�mP�R�&<n�%4�d�e��!��p��Lq8�Ѩd���f=�4U6�م>� q�gKp��)�"�V�+��]���d��@w&ǥ)�}�ѐ�ѿ��6`�|k�E��1>@L�(^��H4d��1qBng�Ή��'�Ig̢ }�jY��LfK�� '��M¬9^��"��7׹k^�w �S[ag�ԝf�A�Į
�ݙN��2�F��	?��$([��P�-�U�fz{=$��&�E��s̜��]N�i�#~��h�$�� �����7l�M�e�n����M�F�+M~o��w������y6��S�-G="Y�=���^'C?��LS$q��M=�����)sf����D�*h��X���m������%s^A�c��.&^S�g*�ִ�G.M�Я,�E��vNe�g�Z8cd}a����]�T=�-���AI�6�����Tq-��3���je�q���t��n�-�4ъ<�UX�{��c�^�����
�l�{�5��4Z��+6���?�CR9�7C���
}��j�@��y[hT����i�����t���i���h�V�Tf&�������V����3�"i���vd\�w����S�O �ۂ�#nN̩Ukc?�8�;���;3��W�h�8�z5Q���}"l���+���d�v���WzP�95�m���D=�.�Nu���n4n�'�g��%7����(�\�k(8���<(��F��}�xbuD���S�X8��􁌵�5���n�2�*���׮���� �"�t�t �9��d/X�B��Elt3��.7��R�85N����6�f�F����r���x���P����y�F��$���?�ןz�f,�7��g�i�yfx{�G0/pZ���2ߚ-�Ʒ�)���C��~�����oA�Sq^��"�R4����{��5~J��l��@����.�wG�u�p'�Űi\a �
�JH�*J�%N�h�y�N���}�A�S��w���!B���u�3��|R�/����AӮS@Ybd�6t_~���n��I[^�9L���'�S-�v�ߖstm��LAE3<
ݜ�eD�<B�v7 mߍ��%���Ђ������>еP"�w�臜�`�Z$VmN�~\�ʟ<�����+J��T[x��-�۲���ׄ>R��a`~l|sfǃ��KYr�c|U��vq�b�����	"S��f@S5/��+�l���)_Қ���je+�eT��٘�z#"ʴ]�� 8߸�����[�A{�J�Z�W���^h�m�K�mmIᾟ�K�A&�R�تs8_T��&+«zi]�ޝ,��E�.�8ye�a�|1��"]�ɮ�3Xљ���U2}�/���=�Tc�����i�lJ��;9��+V��s$<�y��j{�T�D�D����H������`�V�j����\�,X*tg<�������'�>!5A*�M��&?U�Z#n�bU�t@?`"Ȣ���-u'�e��r�D!��`��nL���xּ�l� �S�a���W{�X[�H�l�Ph�%�Kͯ��&s����%L�	RI�<�>�:�@{	�.W�`c�D��p�a5��N-�i���Q��T�w�K�i�S�0S� �T��}���9��`������G�qz��i��9�R��6��rJ���h��0�2[HV�R�wI)��<2q�vL7��K!
��'+êb��C�+�tF��N��|;[ֽ��El��Z���Mb�v�����2�.D����Jߦ��4�p�s|�O��Pu�n�-������!�ۑ*��Oκ���5iZJ�Y�ds�></�C�&��^�?�~���tH�p4�P�[R��_�Y96����T�~�N߳�)��Us��B���HH�x3'���y�E`��g�&�S`Y�4]����=nљ�\S����vh��<�$�}N*��ۭ

��`��x��q2$��(�j�A>�_�]9��>��LIo�C� ��E�:܁y�7���܅�Ā2]>�[>��.e�1���l7��5U>�Y�x	z�_,�0��%��,�����M� (*G9�6n�@��;��T��b3�Ry�h��O����UIgd�lN�0��_�Ro�܎!S�OQɐ����)�
�C����Wџ�fd;���qW�
	��a��?VUJ��'�j]�aW� -���c���{��1�d~h��C'ؙFE}wu"k֋�9�j�i�#��[C���{�r!�ݣ�T��P���\��qʏ������";g���f��Q����%��1��"�<��O8aa�7��s){�+��7W����D��iR��bzo\��9�V��tm�J��|9�[8!jC��
�a�d[>�ӧx�[�jֈ���/�-���s��K(<a,aq�|�>P��L4�I����

F�
P51z�� ����A�E;R����K����D�7�H��[(�-ƶ؋Z���P�`3%�$���N������m�C�)��������?D��_B������6Hh�:8Š(�߂Q���x}�qM7-� ��#�Sr�K�R6�p-Q���ke;~e��|>%Y,f+E�k�l�ּ���{���g~�]�G� 	+��cv�B§0����ty���<���4�d����x���3�}y�g�ЌK�B�2l�On�"����\��������"���'�����활K|e���1܌��~L��΍�k׎��Y�N����7��K�e�{R[���70=ɮ�h[f�͙$��N�q��Ch���?�����X�j��梒���o�Lq	�Q�ݰ�������;�`��d��b�xiN�&%y8��uX�b[8.��	�u�{����=�$��g'��ܵ��$%�-Z9�eN=*�\z:�2#��;dq��X���~̫�xR�'7����B=��K��@B�H�rxR����B�D%�FE��W�Jj�eUt�S��v�Ց�JtΩ���r�Du��+�x��`���k���c	&k)��
�h��y�-/�5�١�,�&Aʬ�G����
ў�8�X(϶��� �vT��i�Php{���\��ݱU0%��e�# ��+��*�9�A�c�C���h��6*۷)��h������p��\�O�XS++a��b\ <w�}�����'kϛϿ
!Di���qzc�Yװn�B^DGU�ܭ��ME�i� ����~�O�`=Q��X����$��MZ��\3,�4o�������?9��/q�2^�F��a�����x�=P}�?���B�ܭ�Z���������[(h?�=l��y�i��|95)��t�4�V���C��M3��P��K�Ԥ#��ݾ��"��&���ӭ㍌>�O��=���x,��]o�j�	�������C�o*��4������,�Sű	���n��ڇ,)���B�Pw�-�CH}##)��jo��;���F����0(o�g�T����������j�q(tn''���SmUͳv��*�Xŧ���%��+r��8�I"`9�Đ�(T�yF��2,�s�+k��w�	{1�˄/��2��j�9(�*�X�p�r���;�'ⲓ��r]I���b��߁���%�]@7��n�--��a�h�7�#yj�~�07�d�ukvA������,���N�ծ� �M�����p9�$P�����c���>�_�ɭ�8\a��Eqjn�8����F688��\ �%ܨtw��vH�int�.��Z\G�@�o�q���QT\m�j�>R�Ң=�W����h
��t�lGh�i���]n�o�^�1���/
~�����1�~��7�݁a�ܤl�E�F/By��s��b��!�1�5���$�2�|o��m�[�!| 2;��0�L��#��[DXȎh{t7'N�2"޿�*>{�Gz�%L�\�xe�Ɏ7��!*{׏l�zk��.��ٴ�ϫ�>����K-�S��ڋ��I;�B�bN,+cp�%�b+zs����i�z�orJ_B6u�̲��']J�h���	[�5 �;9Qh�[Y�#O��b�&|��+�L��Cm����,�w��V���m�艬[��Q����Ф������'��`����2j�̌ˑVvG��a�	�K����;w���~6�V��=4�,D'��9���J�dΒ	�{�"�*��v��8�âd�7w��.�`�<؁B�#3������}O�_v@�@z�R2��(C��o;�Ͻ��\�6~�OX{�)�n����!��7��m瑚~�a�-z� �8�,�M���u���"���c.����������?y�Ѹ��'j%%�+R8�Yv�ʬ���I<|�����{M�~�-be#;bq�cO�'�L����yIɹ��f�$��,���䄒�[��?�J3���,����Sv�s�	6�b�u]N8�\o~)�?�d�p���*є"oi�A#^�.y��	����]4�8��vMIP��,f@M��_�OOc����|��H�n��tʳ�Oy!=U�%Yi�ᕼ򜮳{�+Q�"b���2�I���ʶ�|,[��� �B�����հ�M.��=u.ɣ�"��9XlxVHYEB    4f27     d40�k�6�|�
&�}L�!�ʰ���t,�L�v��;����:�p�X-�:d��D�>�O�B�i*P|NeQ.v�ᖤH�ְ�̓f��О켓�)��Ģ�(S��������Z���T~�����EǼ_=6Gv�Gw���@�f�� 2�ղFs\�ݺZ�3tY[fK����ͩC;0���p�0"�2>|�5�k�������Q��B�3����Mx���e��[�q����RM`_b��s����}]�S#�N(�_ˬ>�mE]�g~���+�� V`wB)�R6����jK����~�l7Q��MZgŔQ�H���W�mp2��xֱ����z[s��'	P)\m��U^qJ��S�4�.�[��BAL��5퐳�׽�+�d@����R����5ތuQ���~	�AW����TP�d���@�f{�"D�� ���Ӄ� �#Ux=D�p�,UX�[�c���Y�^������Ҁ�~����.N��x��l�z�CM�l��7�*��K{�W3.4k+����<l7D~s�h�Lfm�ENj4@�C��W[�'WY7��,K͒����j������:*ku�ªD�����n����Њ���[x�!2ܔ����W�������s��)��nMY~�1,���ƍ>�(�l#\�V���_��̝&q�U�򺵥��-�설d��9�|_+|� �I���V�=S�&�#���(�|�CJ�@ju/SU�F":.�%�$�a7�?�d��H��}B�&�ٝ
�eއ�!�CӲ����>z��q��^)��G����z^[�`3�R LR��<5�W,�T�)O�-@j(��W�hs�IX�L��b�G��)�7�I����2E��������A�d�D�l<�����d.u�TM�2�(:(G���l�n��W�2d����RX:$�f�$D(eF�c��ğ�>�m��C-$CET�\�K|�N�|��7SBy���/�%4.��	*anI��&��I�(N��_�Yq����GC܅ ��K�;���w�+�����*<����Ƈ�0	�#��	!ڦ�X�pݛM-� ���O��ߢ�K
2¾E��σ.QRJ38u/_�����@�\�A%J�G��}��H��r���D�؅��/M�u�:n*:c�����"�p q'ν��c�!QHEv_uTd?�P�'�C��)�|
�̫AӅ!��� Y�5Ǹ�!%�A�{)���*��(Ob�e����O^��lZ��R��*1�ܼ��I
��Cxg^�p��ZP�?+�$���!-�����d��en�U�͈|:���s���D* ��W\��h�}��j��L���͘�<a��LH����F��"����V���YGՌI��n�i-���be�a%~q�dS:dwj��C�j�E֡T�Q�й���M��(�Kzc��s��3��(v[��e1
�^��<�C��G�	3醭3[�X��8S<t��Q��L1�yJcܼٳmD��w͚yXҡ����h��������¨Q�0���cNQ����ȟ;�nO��f�"�?��ٯ�Z��zy�D��ZV�V�,6Z�ڱ�E�H��R���.F:9����ٻ@�7٬���S��?�����8�j��H�:�2i���/8ȿ���N�G'�?6�T�	�Xȁ��xV� �}r�ˆR�������R�B�R�s��?��ۥU��L�n�t�qϹX9�ǚ�������R��
%Hݽ
��E�}l�_�#�F��v���R�>#���y@�	���^[���4�{��y8'~�c.�A���<2��|���}�3�B��}7HS�xQV A��M>�[����K���A#���`�t�wM�;�����8�`u�z,J��9��#w�L��V��W�=9UGV����~ެ]L.{I lyy��ƂI����)Դ/���f0��-~���nS�3���?T>�g���!��hu���2v��������x�2�R/�x� ����3L� �S�AN�k.F�h�jLV�S9��{�C����j�|g�83ւvx�L��c���/}���Z"�"�%��z���y������z̺�\�p����\�:Z���dA:�B��MZw�b������2�>�3�ċ(�D��W0��P�j;K|uP��B� <�),�#%gŢ�1P]"#���ג�.Z��?Y&`��7���J�������3v7|�|���vh3둖�ȋ�"�ׁͯ)1�*�l�U��8Y|�2�k���w������7N����?����W:�T�侇/O���.c�>�業g�>�h�txx,��yA1s��e�� �{6�0�
��o`��U0��:����|.|T4r��נ���*�+>�H�Id��
�F�2�ٮ � �����	�6�_�\��]��N���Q�Ӽ�tM���Μ
������K�ۍ�|q�[YF�z�����%�%dL��ס�B��'Bz����^��������ؿ�
^�@�M�q6�(��mSY��}�rhl#Kn%��B��3�^�\X��N��%�2'�C/�ض�pBc�iA�X���s�VK���Mٮf�)��c�=r\:�@um�?����עzJ��l�r�������{GY�1 	���ul�s�9*&�2����D�l]�34�i��ʛZ��>���#c�}@QLk4�)��1����G^�\���8D�����a�p���f��݈���m�jjS�IV�;��b�T�m{��=�,g� ,�eS,
�� �<��m�T�=t�r?瘐��M1�t�+�\z���-f���e�c��F$�#/F'�"��4��g.����u���Gٓ���Ĺ�'��;�c�+���h���[g���`I�Q��a�b�<����ˡn�:���aɤ�=��{�t3������I�f+2��J�-AcZ?����@=����џ��p�� ���A�1�s�{�*���Iy�J���i�����\�ي��+^�o�+_c�[�l���Z_>Ɋ�>�?�3�Aq���P=�ryԜ+�`���r�,$Lܔ��eZ�7��N��m��ֳ*��F�F��Pc�=C��pٶy�a�9K�YW��#�e��K�� L�i���y$����]D��f�'��O�〓 �§�*�W,�˹ hwś8�`_�cGH=[p%��ء�.�1!,c������F�f�'��P�#b�c�v�#�6��V21�|-<�E?US�|�L^�P#��?�' ^�!fy�&�VԕS�SB���x�{�t�K&7�`	�&�3E���a�}�����ߤ/�oS�?�[7�5p)#��2�CS��� &{��ݸ
B[M;TU��kT����'i&(�t.(