XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��1�a3�A�0����g����f:Ћ:�ɻ	����Z�� v��+�������W{7no�w�Y��-Fs��;Աڈ�w�܋��e~Qa�^�{u�iD�&Q����N�X.s�G}F4�~����9��KW�Φ�@����d�<��6侍�Us�����h�ʅ;]\�υ�d5!������
�K�bLV���p�!��G�S��8*h�
���F���R�Z:��D��]g�_�}NP��G=W��/)�3�����7�����r���kP�[e+�#�|$��HBƋ43[�^ߋ:�p�9�H�ʕ3��-`뻼��~G�0��F��5�e�*�~Q�Yz��ܜI�?����=*=���#d�ׂII���W@��ogZ���h��*�p�n˞8���)Q�y��q.�GH�õb⺂��\�;%��n?�uO�&�K��VI�#��z��q�dK��l",�+��lA��M�V�%ݰlx4XR�dGQ,�,��9r����ٓ����u!��?��7�Ɏ7�l�7cY��#zчS ��f��Y���I⠙(*���z'ݣ8���m5��=����!��ȍ�G�}�0�_����BrY�7 ��l� ��,�^�#�N�Jg�b,��N��gN;�]����b	�"�Vӂ����j~��*����C}<��M�@�X&e�#�7ʹ6�n)#�<K�f,� ���&	,m^g�t�H�9��.�Za�F�Wftq���-��#U�V������Z�
|+��ہ��Vh`�8XlxVHYEB    1427     840
�AH:�H�X�;�xO5��4��N�Bb��Ҍ���H�^F���|v��,$�	m�V��ӓ��~&�I�լ	i��M�pf"�[��7I�'���#J�5���OZo�2R�!�$��Y%���R]����Օ�����%6}x�S��������yҕ�0K
]G;��F�Ъ.�����~��]A��&X��l�.h�-[!����y�9� ��E���|'Tn�K��dF�=�	�������(<�"H�4T��>�3�}GU�'hg�}�CR�K�E����l�x��dW���p"�7�,6�MN���F������dk�{gY5x ���K}�HΟ	#� �>�&�\¯I.B��:/	Go����̗��YF"�4nݭr�NDYU����g�t�e�Y%���>m�#���t�5�� ',�7M�S+Yv��TE�`��	���잊eX�M?��ou�j0D�	�f�!�h.8�T!]�~
���a�<(@�"�u>x�3�n�����T�1� ������;�-
��CW�����UG�cY;��z+�еg X�8����s�������a����T;1�[!U��=��iSY�|z	"u�+�'<��,%k�
��EA��^�=l���|��d7�	
��܀�
�d�j�s�Y���2k��ě���6}�E���M��TW�z����PM�%��UwjԔ�d��g�O���N���%���>]���X�m҃ ����2t����(��Sܠ�k�$y-]�;����Qa�N��t�`h��D�,������ے�A�O.�Xb �����,�fѬF:_�h�*���Hs3�1��;<c4�ܾP�a��ˡ6�%~c.ѩ�f��]q������L�sf�?]�
����a��\C�8��{��޺��5�	�F@k}�_���^d�Ȟ�ށ7��c��0-�r���+?05��G��?����d���BO2H��4�x��=3[~����w�b<�I� s��Zź��w�]�����\	Yٜ9 �8a*�^��Q�`N���n�2!u�\�1���AS��RX�Oy�.��1�/�⩧�7�:�Ln5 �����j!�K���8����*E�ǽ��[�c��x"1��E����0��%��b2v�b�g��Fo�wk-N��;�b�&��꜓)[D��^�8�`�6����)�Q��6�u���<�*vu��*wO 	�f,���|��q����zsXT+L[�>S饔D�F��?c�!w��lP}�-��"��b�҉�A��~ �m���{�pYa���r���a�vl��2�2��塂!�F�i7���HW��j;���}m���zY*�ܯ��B�v�+Ħ��OEН}���1����\o|F|ε04�P�ʻ}ua\
�����d��t׌��꾄Df��ۮP=<�F�G�>DKK���6}׀�.ő���E��hi6���7`3�u��C��](���*���9�{����&;��|D�k��3K�!<�=�[W\��D�)w,�u�^�=g���|�/rN�S���9�U
";��Bң�c��$�7x�*��E��zFD���1���z鮂�N��h�i�lgOYu\� ����Z�zj�XC���`+���c���Y��tu��{���?���p�nΣ��%�ͺ�߈�,X�3I�H������^���D2 м�s=�Y����]��H��;��@�-�C�\�]�j�_��ҿ�W<��O���g�+4(_����W(̙�竆p��EԑM���4���a���>I���ns��.�rh��\�F)w��[B�yC2�yQ+\+R�@�F �3�
���3��QP��shz��Sr��A��0C�B��8��W�xj�
��?�Pu����~s�X�aS4�5On']|��S�3�_�W�_1k="�a�7r4����I����r��-	�ec�&.;6 y�6�0"	~?��V���I��G���EK��dYU�uʑsb5|(��Lڦ��ǯue��<�2�����c�њ��#Q,:�1�C�RO��/��C\`�����