XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��u_���tu�Y�1��n�#Tl��� ���.t��wM���*b�U�yv[ЛE�G�rz���x�xRD�CK\\�2����+L�s Lkۃ����K͢DkU�b���$%���\��̏���k��F�Y�߽��vX[��� Qy�����x}�?gOF�ї�|�V_�}�O��]��M.��T_X�#Uh�� FNa{�����S�n�.������N�HN���'�q�aI��r��X�Ӎ*�u�������	d�0q�Vr��?y3�7�^�1SREߟ�?-B ����@���UZ�'��������37�xg#����!&�ί��
�����oB`-��5�J�3�{����À��|9F��¸��Vr1��� �M�5Au<�LάN
5�i��/@���I1�!���R�ِ����R�?��7��Ձ��Y<�Ck@L1@Զ�d��հ��vD�>��B������^? �*[W���MK�T�G�+7��Ԙ�'��o֪)͌(��ا�i<���h�	�L���:��Āb�$}���B�������n�}�0$��̡֨�'�r���cg��NJ?��ET�L����y-zb!���?��E�^9�g��	�u�;�������M=��W��G��oK ��7�o/G��U����3�-��Z%F)�Qb�{gQY�= <F{�PE�"��-�mO?��ā"��ot(�޷OI�EY���.��T���[�1t���q�Ns���Z��hԑ��� ���N����8QXlxVHYEB    aa31    1e40��]8�daG�]���>��b��:���O]�����y0W�Տɍűd���l9<Pa�'��k��Pv��/�l�s5Fv���lԜp0�/��Y��� �:�|�Ÿ��U)��b���{�#w>J����`��ѻ�P�k3�ވi���V=��kX>�5�d����'*�3�eaA7��h���ֱ}wx0{��6���+�|(a�	)��v
	�� ��QT7�4:�h�ć�T^���7��hU\L^��W`���x����p��P��G�u�(9V�S�.J"$�@I�;*U�!j��Ç�^�{�
��.fMY�XV	7��.u���+.�4p��K�p���$�t�.�|��$�v�y��9ޚ�u6�M��BI�R#2� �	=཰� X�q�b�o��&�,ST���lߚ㩪�e�>�a�+��w$��Tz�����=
2�Fb�o,��^,Ov_Mz�#��� vy"I�{�N�X�{,�Ey��.>���{�XgC�l�f�)��?n�u���m�UO�����l�m�Mk��6�h<�0���0�u~����w w2�j�I�D�@6��Uq��f��'���g�U�m�R�ܑ��U|n�C�8p����_/��s���,]��������}(Ե���ͺY���7�\1������ݣ��/��4�Ju�,�S�˳�fl�a
��ܳj����	��H�A
��Y�%����lYM�[J**��i��i�B�P�B��mV83l4��2E�w'&j.�hk3�rͶ��7gA�C����I��b��b�����9�bJ5߈��:���{����=2T�=)�C�T~w���x1I�����+l��W�A��\�J�6�!�z��p˨�Ȱ�AΛ�8�W�_E��>��^ v1G `�ӽ�t���{��Z�XT:�
�AA:Pҋav�	�ʪ_���ebǛ�U'�[%�Oj�a1�R2^C�<��ԍ��!oA/��^g!O���]��G���i�;�_;Z�	�!/��]�L
�;r��N*+��8^Ћ׭N[�Pn;�-��?'z�P�e񥂒H�Cب�?��*�ƭ����H�
�w��XL����yN�Ñ̾W.P|��<���g�;hO� P���Y�E:?{�!�]K�^�ٚ�@ꯙ�&��\���3�J���E%���0Q�7a�F[\R��xxp�|����~��?�N+����ò��I&bQ۴d�0�|-�L�o��1�U�w��Qp�������\���Q�N��U���`���0vv������)��d�;nߌo|]I�C6{�(\�q�XN�#��!�	R̖����I坋�aO�:�7u��r?�K�
��-OMcD�%�6{
D>�H@;��|cC������[�2M����5�=�L��"݅��0����5Y��g�p1�:: ���#m��F���K M�K��Za��s)�U�|UG�?dD<��ܩ.;��)�su@�؞��4ڱ�3��䙫N}�>�.w��h5�J>��B��1�ws�R�F�0�����ھ*�Ӡ~�z �����mO�ڐ/�P�h RF�h�(9҃|��-Or�|+�����p�,a�8�i&Ϲm��uj`zr�3I��-���]���������g�����	�
��DZ�n�O!������Za�e�iˑ��JL%��j���QnW\}#�Nj�B�����=��?�qKFS�C�e!U�'�m�x09���K�k��&���6�@�+yF�+�*��ѣ!CdO���A#�w������^>����Zً�WnG�n)̥�i\�K]��w'0�[
$��/��T���T�y庌���]@{\��3���j+��ݰ�����f�D�9�Q�= {�}� ���mC�6ӌ}3���&����C���5tC��T�q�|�0�4�gի"��'����_�c��/Ĵ?a`lK��=����{���E���j�@M�*HMI���! =��.�l��Bm���IߙԈ֫��U�H8=q��G��� ńH2�b�Mt����9�ke�z:�³@˱�T��CIRV&B|T��TEc�gl�K���ٻ��~5���k�5Q��g#�u������5�si������C���K?�"׹Hε�'��~�չ�ITf��hg����%����k/�~��?���,�(����l���aT-��1β ��Hj���T.��w��H���Sz�xM���K&�9 s�c��%���(G�o�^��9UE���]?ԥ�n���\ͨ�Ի�H&P��[�&��wd�m��Z�B���u�e!��HF�W"�R񴜓*��;{Jh
��!=�jsm//ѝ ޜ��@E�
Q��ɤB��#�B���;��aV!�IU�BW���;Ч=��gǪ��C�%٣�v�1E�)�O�x������Iq���CT��$�wc|�kE�6&p�3��*(�>�����-d#�1���ʀ�	���q��,9����|P���)�͎Y�n۲�]�DJ`1� xWs�gp��F�$ǩ)�2s&j"'Ď�d4��,:���������Y�NI����ߟ����2���%�M��.�>'����u��[L����2l�K�^vq_7�JT/��&�$T_GX�'wS�&���~��XA�oK;S�S�-�'đ�~~����zXX�d���ȟ��]%�������~������S=D/���S%�fR���d����]6KD�fz߹��.؈�.��T�Q��rܠ�Z��D��4Bl����������=��1����+	%�E��[ߎ|F9da��eBD)�#[)�tV�~���e�v���]��;�Zl(%�~.�k8	.W�Z��@ff�~����Zk�FQ��H�8���Y��E�X��" E	4_��riS0��{�<Pv�p�o�9�Z��������*@j����ԗ(FR�̴���q�¦/l�{�沃���H�ц&v�<�:5�Lg6Zu�[H��`)�6`{�rBp��r���/�ݐ�Pb{46�=pW��J5������V3=��$D`�UU�u]l$������P~��%EW�$�=�ˣA��G8��ϕfof%]�"��!�)���Uo�P��K�R;!�L28��i�� U w/c��n���#d��y粍��aO�%���~)��zj�|�	�I���6�X�N_��7��$:[w#���%[�9��<���ɼ���\� 9���M�a�2�N�7.0����d��X��R��ow�<��n��Q����B� Q҂�~	NG�o�jW"RJ������k�2���E�ڭ���|~2�D�+��-ۆ<��+�w����"���h��)�����7�8Cc'wPe�o{���wl����Y_���<b�����	O؞.ġy-�И>���W5��!]Z�jBA
�1S��»Z.�X���U�,�!��1�C���vE�@6��[s�g��N�v�g�}T�
!�ds�ew�Y�N0B��u'�/ ���bC�l�O�f�^=Pr�QxPv�[����o%fc|�����Ъ}����<ln^I��ܝBF�U�x�_���*3*�%�/�P���w�SYVI�"G�}����]��]���#���$A�/F@�$I,f�c���4�~�p~~X�vI�BS)���\�Q7vp���4�kY��;؇����� �
D�+R����u�k�]���D�u^�=E�y~r�Q^>L��LO��Q<������5&�(�b  ���NP���-d��h��.����ʌ�K��ե
�B6l�1��?P�Wd|�/^|"�7Ϣ���'�AQe�����IA���B�b�d._��"�s��p^~�]�]�IZh�����X�n�<�Hi}�w�}o�cj���$_�;��!��$�R��1z1��}kI�L����*�XFE��
G��*�i��o�X�)X�l�t��)��a�j:�Y���Z�hU�1�v�.j�a�*��*8Վ�z��ta�F����t�Sۧ�ࣇ��ƨ�2o5� ոIXq#U0`m6~W2�!�@��C�B��ؗ1u:��!v�X`F^q}x(io��1���2]� �~a�Rfѓ��Q�!
M�i˩���y�'5�R���o�B���hw,�!�ş�UX��V�3��b��7"*�c�kȳx�C�y�v1	F���5������%��Yd@}�&���ӆ�&)�;xl~S|���^�;8�Q<{ <���S�0�^���'����l�E�i��J7ͳ������?�����_�&�=Ac\�{����w8J���k��B��G̅��y�����/eǙ_VGo��=�u�a����_�$�ӐG�%�YO����R�4��kqQQ�Dڭ?a����G�={��uS}�n��R�R�T f����"-�Wz�2֒n�;���v�?%[����]v<&�6��+�@^Ѹ�>gt1\R�͉GǏ��c�˂��e_��؀ཽ3З�0�M	�O:�+�+�h
{u�s�0�G�M��5<�
w����L��s2N���c��E{c<��p��rJ���׭����H���BJ���
���z�nd�շu��-���` �}�ߒO_�<M��}��ld�^#B�C4)tRGQ5]��~�>[�Ĩ&5ެ�L�'���ͪz�(�0��m����[d��2pN�8x�C'C�C��N(�;\��l��n�L�� jF����5JYbf/� ��9��T�R~��(��x2J#�&�U��p(+Ct��v�3'�����l���5\����@� �̡ͣ�^��q/�+�+����)��YCZ�K^2����{��_0c؎X*�o�43r&��H�IL�������b�X���O��ag�����.��N=:���	��.�~�[���+����lUD��$Ar�?�&9ؖ���1E��`�]�?�I�E� 8BR[�Փ�m���%�"�G�_rV��JY�ۉ�L;��E����(,�O��<�pS�
u�0%�0�f�X�����"L�mO[h<qU��wzO@:��Ca}SU48�*�8�C*�5d�ӈ�O!��VT�l� �qCTNS�wRE��~������΢�t�̘c��4j=�6��5Rð]���a�]`cq
�|����� ��9*����ԣqכe��YB��Q��0�1y[ �;0n�6��!�T�G��p�W�XH	S�Y�:%,���PE���md9�\�6x��}b]��������=C�n=�T��rvD��wT��2f�W΂U�D�R���	X���)I��^!����o4����Gа6J\���/OQ�TJ��0;��ɓ�����\C���Ԡ�h�q�6��.��������;�P�=�y1:�Θ:�L��]J�\)r��^M�^����.u��i%!�Q��]�.:FY��HсW�,� %,�E?��z<���",J���YcQ֫P:�I��F�R�[����|�n�Dx�x%zBa@�)��0�d'�e���`
���;T�]�s�X�~����D�zX�x<A"�]�������\Nv���X���Be�_�㜴�k8�����X[���S�%��ӌ��N:�ߊA��I{`좗�8�Y���(t�?c����$���QLP�����g˒��AY�1xCD����]Uތ�����("r۶��7�ޖxe ��'�n��@��S�Y��j��� �k�6c�ث�:���t�j�rS[Tֆ�����M�F�0%v*� O+<����a�=����|T�t�^��0�iD���a���L���šg���x��q��C(��*���|~��.��Z������3�4]T~� r!�%�3�]ߌ�;��V(�V�sa��C�(LؼF��rٞ�������dMѪ����TO��tH��O�J�W
�׈}�Q0�����M���r*���p
� E�u�Y�.����"�H��U>V�Ҡ��P�q^�=�I2\�G}A��'���ۆ��M6�|>	��+�����F;�����<a�Iج�������I�;z��B�#��A%�^�D��ݖY� 7��Q��n�{qCIG�ȧi®�]���lº{��@'��>�4byj��3Mv��3�hss)rL���#:�w��0��;=�4O8�COo��BЇb8.Q�[��Ejc��o����W�s~0�n�yb�*~���:D�*�pb�qc�(��$A���C�g���$�-O��hΜ^�z��eN�K�B��
Û"���')��"h۳���eC=�E���U����]�81k��6�����Ӡ���� �&�xb�n�9A��|��8�Wc��5ڠ9;�I�]R�Zb������ڟ\��Ⱦ^4�s�-�>����H�`���M�oMR�m;��u}/<v��Zɵ��sT9��з�J��:��������C�31�l�̢�昜�$OL瘋�a��)�Jf���cQlyQN����W��X�]��R`f�k�ʌ��0�BY��ے҇��з|��8�C#�B�M��I�+�#֨-�<��2�E��TS!i��o�1<bk�م\�Z-�����")���$<>�����J�>
q�Ԫc�Q�3ɾ�a�^-��|y�רb��o�Cv�4��BN��F�"�j�J�e����xڒ�t�ږ��|�����B�&�����z������������`#���GW/�>�T����5E
k����BL1�r�ū����X[���0�v��k�3������=������A"�#)l�=H,���I*��,\1<Gȹw�A �`x
#A]h~E�<���R}u��׫�.h�&~��;�Q�IM�_K��J��g#���������)��6����7G��l��58�����ݭ����2G�K�{W��d(�5�K�[�)�!������mz#�`�����G�Tgs�>"/$��#��V��cW��nctG]�����#3Z\td	#`MU����)�F�4�Z�|r���H�kB�i��c�;������h��C
,�8N���I�3�D�:䙸ς��'�uJ��t�RQ�ӊ馭u �dP9Q:ހ����<�;a�����-E/rMԺl=��H��r���a�z��9B^~�d�b�Xl�wצ�Ɍ��a�����5'U��`�N9�� �~v��gT�H+�!t=ɍ��bm����r��/�%dt�S�p�"�_��22E���c�v�#�F����nB�@.�(A���T,e���Y`�:�bbf��f)����p�3|��xm�Qr�k
 df�� ���	�;�H� ��z�0�GM��P�����z1��$<7��-� H�5���p��T�9=�*dp�J3ڼ3�Ǥ	�rS�%���@�%{��b�l���J�C�.a�P��v���P�x��eĩ\2����s�s 	�O�K��r`p�

�<����Y��4���:q�QgX�t"�2���@]4ɞ��:P��'��`�r��<s�u��e��w*���/Oa��� �Ɉ��t���d#N1�������6X��ܑO�B鉮��LԀʜM��Q��< �4����*�~biF-ڽ