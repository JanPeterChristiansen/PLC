XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/�#�y�Mǳ���i�@$Z�Fz���ϲ�e@51�:�s��Q�Ǘ�f�ye��̴���q�Y����8�c�~��x�����՜�v�:�x�J"��hҲ#���G&&��3$q���r�yή�IxoV_�̘���D-[[�>�譝�N������t�u�Q��>�p.3��(��ޭW9@�)���N����u8wJ���5軆�A4�~�W�]]��Bq^��m�:�l��
�	�Z�Թ�
���U�gسp;;�*?fTm����J��Ck7#�ln���U�$ݺ *#�(A�U'�m���GS
�j�P�{�ũ�,��,�}�Ba�Ng��Ε:�D\�:)x�~	dU!���5�Gl��Z'�{SFD�1?8���#7������u(����$���dcִ9��4��?���K��|���ϕ�y��|)%�6@t�j3�6���+���m�Iǽ�`,�]"Z�H��|"�e������e��q�r��o7 k'⿺zUPsv-��&�Aj
i\�Y%5)�ܒa�1<��OJ�N�ډB�:F�?XGX6��OXq��K�DC�ü���>��"'��@���B>M7�u,�E[����d8hCL9;���F���R����!D�&9�e�":��s!�G�B�1�0����C�FݹC`�C��h'f��ă�t��=[,�U���U�n�7�'�;�q�eGo9��4G���ȓ�W0�;vnS�L<���a�a�x1}s�g8w��0g��~XlxVHYEB    fa00    2480{�C$ �;;8�~�`a3ٙQ�(�D���F;y��qR�X
6)3�Sk���8ՃU-Q=�MuL�J��q;*'�͒���S#�U�����
�T�`�A�
aZ7��a-�W'6l�ƛ>�������MV���i�SW��ZA�:(��Tg��W��5c�4JŁ��oU�D2�S���@b�)�	F ��^�
WyVOl��mu\�X���X#Ň*�N���C�Y__Ey�H�Ȅ�O6�ђ�R�.�w��Ug�LN����%��l�\`��o�������dn Ð�<��tδ�))y}�b:���X����o?��Hh��q�'�%�C%.���! " �E��gג��p��܀��XW�\����F��(�*�$����$��/ F��!�W��IA��#IsfmPkGq��h	����·�˖n	�uL�GYUq��!��b1�"�~�;2�4��7��q���TX^܂U$�f���s�\��n&*�dJG
L�N6ij����􉯜a^��n,$G�?،��K7t�6��6����m�h�5��&�X���_;+W�!��;��p����aw�nm�B�#)��>�Q�x���\��*W�<�DN���^�=-C���}h�|��e.I�K�"[��Q���>f����M���dAwR�0%￙i��x����z�Ā��j."	s������&�=�����ǡ��̒J:��6 �	��̶enӹ�TN��S�+�z�����BP֏�	�]2�
!uhu�����j�$ϼ�_��JgD�j�/ �X'w��3��%+��C��w���$�#����X�(���v�,5�Qs�W*;À98n;����~��9�٧� ��[��f�p"D��b�jH�qӗ��0�Jo
�� �ю��+O��k�
{VE�*x�������vq���M	,X�M�y�!5p���A��{�&�"��V���W��iF����4��U�j�a��ǳ,�'��A�oj��.����;���M%�K��2.5N��>,6�w����	�Tk���O��f��GTܳ��t��
�>��O���T~l������j@�'�6�;��7
  x@EG�/�	e��R�r���^TM�"u�=�Y͝�q���M>�^��g4��0��+�
~���AD�����`<���PZ�?hTv?�`�O������GQ���d؀��n�{,������=�z��x�7��M�B�B�n)?]
h��Z�y>B������7n��
pV��/���b���%�u�T\Iۮ��������o�-���Ԣ�q���3�*���6e�Tl�I,>��_��v{�	�]#Hf��qj";>�sa�:��C��p�*���X��b0D�$Zj��޲Ѻ�9P��8�?X_LizL�:L�u�v���ޢrMkC�v,`�� ���D��朂̱⢶.���;v�+�S
��Paশ�3���v�A�!�
�{r�'�/?����=��Zu��9����'j�N��n������G�|�-�ᣏ�-F�����xT�ή(�� �]]Rʈ\�	����s�.�53Һs�hpU-y��$�Zn�c�u�+��Q��HiQ%�h�	�B/�;=v�Σ��隔�i�y)�CpN���3]����o�
���`D���� �UM�]��5-V�-k��Ԭ~Y�3l�Ύ�ޯ?.�'�?ED/n^�@�kcc������y�U�rY��E��;�0�k��#ޑ�������}J�K��]m�'�}��`�տ��j�$�TI:���E��D��]�5B�8�����O�5�.@�0ذ8�a���y!��J�`'g.�F���q��
��f����]v���@$,����C8=4f�Bd$,�)
���\��_���=��� 2X#e7IU��t�Í�-*|�ަ��L�޽�MlQy5�4�!\�h+�l��G';��[mţd�f����l��ϬhD��Ճ.�sO�E-��cRSWB'�G�]��FF����|�૚�����S�ւ�h�pV���c1��G":��Z�A�;YO���M���]���z��D���zv�LPGvF]� ��ɦSJ)�}�(.��{��1���:��F.�0�
�p�^�ݩ��Ѣi?Z@����`�?S΢�_��15��H�;B��f&����͏ �$h�4]@���~t�?�`9�G��k��!9S�;���E���~��Z�5�a��_#� vUD�)
	�h�e�9픜J���U�ۄ���'%����}��ï���`��;��Ra�@�c-�T��!��J�æ�����<���Մ�uK&�+>N�o/��������A��F"SV΀D�/��I6݉�˕i#�����2o���7�1u^��Qţ�z�m9.�|�?�]֠�~�%��p���6orGy��N5�٦�l����6[3�A�8������pJ��3���������m��VS��eΙ�h�1�[��ۨ��j��HP�ܝ?����3^./FG�K�A�)�!hf�ӱ`��lu�X�y/��wvuEG�yP�(��~]|ھ�^̶]:�լO�YM47����M��Y\�d"�DAg�O���`/J�Ɏ�_<b��Ş�f����T��9u)F��b�
Ds	6̧�tc����u�4���5c��i4�3�&}&{�����92��S�Y�D��Rk��,�n��9H�}�V:�u��y)�$��8�xW##s�1�C�����f%tr�
�(Z��BA2$d:+��t&DX�}%o��V=��	íG,��)-h����{n,�~o�D���uP�aiM �;RYY�0��s|����L�GU VU���u獥#�Ћ<l���~��y�j�>���)߱���)�yAckD��X$v>��?��e�ekg��@G��V� cb��'�������N�P[���2�*��mOrY�1fI�.��.�.*,�PN�ݜI�V>0��j6�������E��m�>Ք�a�����.�ԧu����� ��)�����J����Q�y��T,����؊GWO�)�`no�4��#���OIxZ�W�Ңq�R�l�2�h��V�n=J�yD���·Q�$DPD1���	��;0�\E�CaDI��>j��{"<>�Ǯ%�]�\�%7��P;���� ��>��~�5��6wW�3���%s���%6�U��{=F?x�v����^��ZF	�������q��'v��.%$��/*�������C�(�Gؓ�i��4�`u�p�:��ֹ\V95�N9H�!�Gx��ǂ��zݗ�(������4	�1�s�ዿ��Q^�4��B���Ac�՜FX�g@�\ә�-�&M*5C���;�r�^����y�������QU�*m�D�r�1������j4N����x�`E9���#���6�����L���}4�i�]�<DN��%���b��V��)�H����������ʃ�!��QҘ�m/(�#y��t:����:.�N^���j	_[���9���+���*��Z��y}�ϔ�6���=��*�k�g��D�/�>��
����X/�"���)���W�
Q�7�GN��o�W`�Xk}@�~s�ʼ�mPآ᤬ʵY�����x�́��f�J��W�
�]
y�X-���)qd��V���qo�Ty���C�c�]m��N�+�I�LԔ�*}�;�)�RV~p�5dgt�RJC3�.��]f`����^���-_��L����	_��Y��F��]�s��+/&�l2���78��1���D�����k����g�����-��~7c4? ڲ����9!j~P���xP��a9����������SŵƼk�}�����!9c_ʀ�-�q[fÎ��G��e}?y�S��8��*��N�4����;2M(��O_Ʋ���c�޶����d�%����U찆-�j�屧xe�t�J��G6O�}�تp�Y5�ATQ�.r�H]]o�����vrՑ<=�.r�pO)��~��(&,2����%�U��g҉���+ h��[���.�i��� h�K��`z�*��n�.&��uC��t"ׅ��X"cZ��j��I8���ں�440��/�st��^D�%�@��M����mIt����R��Q�:�;
OM�K�0�k+>���-A����&�J6��V��'��;O1
��F��g�l��݇�񚲺�.R�,BM%�C|�%Z~��/��3xQ�Q��#m������
Z���Vz��등�Xήz��^��3��J�$S
���n0�ڋ�x$�i�T!T��B=Ϫ��:�w!\ �������Q(c���"��^%I�j��\Ӗ�虆�=�)O��~�Y��TG�Hn���C9`�D�F h�8g����� kd���h6�>��*�K�(�)c@��R�Đ�fl�Kd/̠23����v�V��I����@b5� ��D�}�3�03.U2�Y��RB�M>�ɽƩ�A�p���c�-�|
�莬B��R��7�6���^���D�iA��I N$�0I0�M���pl�/=��)�y�W���v���H%j���|� ����#�L'�� 1}�ңD�59���MPv�����ע���ʰ&e�+(<̘/�l0�`A<{
�]Ԯ�ˑ�!�RxC��B-h[bh^�gM�X�����T����q��f+��d��R��x����ڑWX�NOu���3��/=۸�����kp�i�$Ng�T5���Y_V�[����  �ۿe��G@�m���ui������z�_dQ4��v�X�E_���+7vP8[��](�z�'�힐JW��Kk��Dr�Gm�Cfsz��I�j�������V\�b�U\3:�ʳ)�\<�MSN=�V��
�tc�<�[�q�Z��c�X^iE�Qc](�ȳ��"I>j�h�D�������-V�Ь@![P~�@9��)���.�2�C����׺97F�}���\�����zx�N�Y���)�f�3�]uG�MR@�3F�e�R�G��ڳãk��~ �2�a�}5<���S��VO)�-���)��ծdKi�c���D[�ܯ�e�m��p��*+�q��/^EB��W/��4�+'���N���8�4����<�� �޺�4�js�+&�D�JD���G*#V�a���{2OP�E��z�a/O����z'Cdx�CM����C|	N���-x�Ϲ)0���)"�z}�aS2�X�"2p�n����K.�ğ�!���N�������P������"��c<)�\�/H��k��N�ka��N:$�z���K�$dBh�����-��KC�t$ݰ�SN���t�������pS�w&B�-[Gߔ�^<l��6 e�^�il��q���=��m�l�?�	��j�J�u��XY����v��$�!�hB��RՀ��o4n��1�� k�S��;�Z�HQ���(�}~X1��2)ֱ?,u�Q��� �ĎD��Q�jC8��)�3�z
���X�mV�$Li'��	�b��m�o� ����h�{r$8v `2!�����%�}��oy��A�_�R�P% ���H����~�S��O;1�5��/����#�DK���'�5|��3_3E��A)G���p�C3$�+�C�-��Չ��HS�W�Oɫe��:�m���w^R	�DiV�#'s0� 9W�aWx�~�����y�Oa[�����jɮЃ��LN�fu�_�Sݨ��#Ku��z��T��i��$y���S�ЍYp҅�-�VU�]�D%��9 ����ƄB<:�k.YT����;�)U�VՕ��}_�׆;�me/�U3�AQ�,ѽ��of�D[����Zo�� J��y}�e�$�����f�&�W#[�$�GK�y3�O��KR6���D��V�&��!����I>��Wr��!0�#�W<)-�RKbt\�$�32�vv�t�!3E���T%��)`�q��R ��\:��HT�x�"_	���GB�"^!�������h����Sւ���q�3/E���wU�C�x���d��ty$�� n��,2�#����N�Y\Fļq屶�Ǩ5�N�(��;z�n����Ǻj�\%}�[Ee=�e�uAi���='�$Q@% ����LͼSF�5}��q��ǌ%r;�ߕ��%(8yMو���l�O��y��1v�Kxc�zi���R�4DOjK�.n.�o.j���!t�(�̼��9��߰3�_��j��� �,��w��hr�˭���U,܆x'g'ίz���,������i���.!�II%�ڻү�N�[�i-��E���R-Ex���C_�t�"P(2L��B��'��OU�va�}}k�ɛ���m�b��+����]��-kX��߰�x/t<�F��t�K�Ȏ��
L�}ԉ��:�H�^ۑ�	mo�K��b�ڟUp%�~�$��ϡ4�,��;�DJ�\M�~E����A��1�H}Z|�W�G�l�	� "����~6�����SA6�4#*FQ�37mz(eLlx���<�\~88�)Ăi	���<(l��˚m��`#����D�Nܖ�����$�)t>�Z����������pYY��2�]S�]��v�humW�I��͗AԠ[�I �9��Zlb� |��H#�y#ER�=�+��K"`c�hݐ~,�����_�y|��3�j?��8%q��φe��+f�����~~F,��<+�6F�+��m>Q]aΒ7S���^wٓ髳���*��zڵ`ά�^ߓ��xTײ	�my��h�	ŵ���
�#`H�����P���|�Jx6��k%Y��.aLնFʞP��C�]|&����E��j(�r*:���1~ޏ�(�E��:�n'��+�<��U���Z�Oa�m���G��K�{�;D�ϗk,rP�m�����ʾ�����R�`��[v{ f�0Pr����((u��+JX19�Z����T�6I&�v�[ҠHB���6�s�(A|uT��躉���v��j���9�y�Y�.XD��A��8>���� Ӝ�՛>A]F3�/�gMi!�E��`���X����P6K��`�V'�>X��L�t�V �q`&�X#��B̓EX=���������ᱳ�9f��hľ>�U$��GBQ;d�bUXw��9\������)B��qp]E�����&ʄ>(O��4�8�:�������x����d�P��ů�\p�-s/\ (Ѷ�#��tQ�cB��:g���zQ��GQ_|���p��x�5c��Nu!�s�s"~�_�F�p�{�g�b�V�%&yp�
Y��u�2����ov7��NL{V�P�#��Z�Ow�t�)?��_��5�V[�lRY� ��s�W���y��T�J\m��8+�K��!Q[ٳFh��a��B.�ރ�� �0�5��M团c�C��\�Q��B��&��|f$y�Sە�}-�xY��s�
z��z����^Pjyo�2��^W�������V��_�#���k�����~�h��"���పcpT�[�cN��u*��[�k�r�&����ƙ�])�bȅmM-8:��Ov�M-ĝn���'Ǉ�n/2h�#�Q��� u`N����Zszѵ�E��_����j5sp����C�l�n��[WT���q��P\�tx�>�oHc�ƪ��M5W\Z���Ҩ��*V'����{_@I�џ�_B��%�v�u��÷���Z><"n4k�*٠sTe��c��'����6�>Ȫ4!,'���t̻a+�ug(d4�G��K%�ɽ8���ޖ���9.���D�J�ӑª"�E�3zt�e��w�蹍�ع�.)`K��T�,"_��{�ج���G��g���%ŮJ��x�(5�O)�h
{���c�H��@�ߨ���݊ڧ�gF�*C��
>��5X��	 ���="��dÎcz����xY�
��:��1�/�0.��wK`��@t�ý�dV��P�k����h�'Z0���͒`�SR2� �W���ܧ��	��7���6����f��z�@�9���_c?�n��2r�xW�=;���˵�3p�7��1�����*T���C���� �yw,*Z�^P(��Z^�߭ �BB�⩷#Q{ڗ�(uR@Ë�n'���1'�3
��R~�����~����󀿙T�4��mGT��M���L�v�f�+��ܛ�y�?�W��㰩�ئ���n�[�+&�G[~+��`��crwr�(J�N�^�v��:��"*x9��G�.f��m
��	�%�ǎ�B�ef�y�U%�7�[{��[%U����� �|
t�^=�[d��{�R-Ao�8��E�]wef�����:@�C��6���'�~��Bm*�U���ܞᒻ�GC�2����B>Ddd`�Y��J��|g`�Q��%���F�]��ڑ�MA�1���v�р4Hp�pd�����qw�z���7����6�B%'�&E$����3v�H��N�9�5ދ���lf�[A@ٸE��|��BeK����$�S����c����)������ft��U���^��OM�3�E���󴡿�"A �6������N1wr �fpu%C���vOG�n*�=�[C��kT�KB���&�$�w�|��I��յ��Cն\�}���fSw}�x�J����p� �*��ʎ��)�J�#H'�2�8#��3�(#0�w*e�%<k`�]s�--r5N��8G�x�R��n|��w�Ld��J5/�S�ϋD�p�i���xhob�{��P�� ������#�7\�B�M-��;��&0���Vq��8t0�� ���,�*����o�0u���Z$*��G�	>���!O�����@oC/�1�X�c��;̢M�q���g���z�k�Uf�(^ʌ�L�e��6ܑF����b�������������^PI�ҙ�糁*���Q�
L�#���wk��9o�z���g��l�c���A���o��%����Y�%�%�6��-9tZ�>蓖�A0�Y��/&=2���9������I���*�buV|弧�a��_�M��e���Nw�0��J�;�8eK��T�=��'��bfY���(�����I-����:�bX�����t���=�{�ˏ�P����Qӂ����x.�XlxVHYEB    964e    1150&�s�W��^v����>��c��.��� ���:Is�����(#kE��Ұ���e�FL\���o����ω�̉����m����Z:�럏qp9��K�u��eZ�$��P 4�5���b�a��>y���鈲[5h2X#���)�����A���W�n)��D�34qQڣ����$i^{`ʠW�Yf�B�Q��PO~��as�X:6/��@��eaeW\py�����m�Ywt��VS�(�.l�+����]Ğ�L�a�8N�@��6�U�����
D�+E��h�x�:o�!;;���o|
	x��R��D4�)ɯ���@��J_HI�=�Ϋr�	`�?|I�c��e��֋�-�V��-u�P��M����/s�6�s�B�c)��3�h�w�Z;����r��I���b��g���%�:�t|��a:����2�x�wY�".�u�܇�Wt��^��W0Z���P�+�Y����!�C���;�d��^�ˎ5�5�`b�e\����&i�E'�Տ��U|dGN��,�8��:��>����<4@B�(nGB�Q���U�H!����(F�ɕ�6'@�Ѩ�j�#*0�v4�;w�a���_���h���=��'�г6U!Qo�L��r���v�����u~N1��PC(<b)��"7 /��F̰UX��6�~l>��u��r@����MPX���7v��81��"ގ	���5-��~P�HR{�b��- J��̃L��BqH��ne�2�.�~b
U2~'�� ��<�˺�k�;�^�Ӣ#{l8�fj�!V����
�}`,:����+�pO}:u��<��[ �)�����#Q�h+Y��r/�Q+
s��%�j`��Z�|Y#jA5>�9-qG�@_ǟ�,(�)��ߢ��v0t�� �-�G����ػ^��@�D�e9ۚ��f��c�_´��g�r/���43>���H\[T�'(��&T�6'�al90�_���p���J7(Ѯ�
��6�y�0��M3:w*���v���B���xi!�j�$�}���W���K9�ZP}�FK؟��fĬ�.Ϋf����O(F|L�~[>�:�93��4��,�_��GFB�+�a������{�� ����B���a�d�^_��Tq��O�!6Y�q1�SL���7��m��Mk���iI����x�O�DW5D$pE�7�o�6�y�iV�>R�%�X�Y���{^�4�~��RJ=�ҙ.2]��+H �D��bBطS�G	7�I2�ӄ~�`��F������a�|T�;<�Av�{��>N/c�U�/)�1�4QA�ስѓ㽟�#.����.u����q�etŬ_G���d�h���>c��pw���1��3��On6#��wq�wt�^r�:Z�x0ֹ�0�K�5�v���3�-��Z��d����pW��J7*��&h@�NXa�D�`ilZ� ��5��d̒M���
$D�y�P�a~S�)BE��rQ�p�~�E���.(ik�Wi��H�K��e��\2y�j���͢BdvC²b�H|��-1҆҄�m����"�v��SS��9ycE�nm�D���Ԭ���9�n���l=֠��2aU���t��p/Iλ��n��Mk�Mʵ�=ҥ��<�´�5zp��b��I�����2���}<��D޲�I��ܥ0��j�5w�/"�c�����k�ԮT5�2�==�3��ڋa�v�wy!D������&p�ùk׏ ����#n�sI#�n,l���pr1����<"�TDcH_�f�#�E��hy0?]��\���MOi$��$f���k-y��ɜsH ��w��	�aB�{c���y)$�w��p��^���zp� ơ�aD�J:p�P�Ul|��V6k.�=ߞ�����OV�O� D���*x��Ցq�zHnӷ�YC.cN鿷*L��42����\�C�E# �w)�Qb;����A���'gF@��ηdla2m��������T8�J��ĄF{g��O��&�5 ��5�S�U��Y�* u|%]BK;"���X�dV�JD��`=���N����`�2|��?�_HF8�s�!��]Ul+���IE�v臞���3�3}�w8�l�:������3��,D~�G�T�G����e}$A�_�n��L��҂b]��'���F�ԝ�_�)	���Mx ==0�����2x�3"�6b<߾3��UR���*� 79��F�� �u>p�HcL�P?��jp�c���������M�+r���i�M��'��~|�*�X����<���c��yzmZ٥񬮓151�ʴ���d�i0νB��nP��`�s���q�Pj){WT `e��Rs$��q\�6f�x��R���^ۏZ[����8��~�s-�Dq?uMP���
��b"!EZf��֋���oz����e�-��M�*�����Ք��:�Ji
�Yd�i�7nꈤ�q'��M&��2�oe� �=�ћs>6��dn*��.����w�8.!���[}0/4�>��D{��Ԭ�z!�H��ɏ�eG���Al���<���q��	ߝlXEG�=�ݣ���-qX�������e�~%ILS�r�p�c�YFj��:�w����r�w�6��eg򞭬�^.���m��K����ȩԪ�Q�������NK��KY���^�4[*mÚ�Td���)r���s(�ª�e39"�1O�`<�F�(�sK_�T�����;�(��8r��a�?Go�ye�M��N�}` z��19�b'k�>��̾)N��N��s �y�1H�K4*�[��ѱu
�9�7%�@��tf�J��R_��V��r��Hz!T1U!���
���I�>;��u��U�wY��Fl��s�6��v=f�ojCu᳞+�!̳�J!a�i8�
�S��'��w�(a&�e���!���*h�2�)��^�z�p�~�="�����F�R���9Աg���bN����[��ލ�j����?Mr6�pfcN���'�yM�fU���66>"��<C�2F�A��rJd�Ě
���܊B���F��bC��,ً�/|�� �y *N���=�G)L!Y�d_]0(��l �F�W]����Q^�u��ףI�˼2��lڈ��8]�}�m�G���?�g�b�����833&P�G�����A,��B���<��5�������꽯���[Ҡ2�-	��2�@P�vb������{�O������Ot����)�����<��OB���Nk\-��܈�ٴ�!��±�L^�H{��s�	�&�rK�xI*��e�pbA.����U�Y�\��� ��{!����{붎���@�Q���˥$�:Wh�k�(�b(|��\4���=�z4��jY���-�X����
�ß.4��Ԯ8jS�{�մ����K݆qF)^�rm��X0�(������z�� E�%�"�+@�c�B��_���:�܆JY>B�&)�~�h�-����{�'G�i�ٗ�TSc�팆J��-��127�eu�d��:���6���^����fWW��T�{�O.#�s!PG���L�Qj�3��К	��d�
8~�-v��lyD.k!��(�'?=&y���J
PE�P�f8�8�����3{��(�=�G�]Rp�'��JO����Jg�ީ�tG���V� r)+���X�>Y��6-�E��:'����Ԛ|p���=�a"���T���.~������o��|z��s/�����}�4�98���n
������͡�鯆��rM��ʇ�)�d���ek�^��c�!/���,�e�+S#��~Q�ٕH\Y��ۓ}��CA�JO!�m�@����1���W[K�xD�ɪmE��N�,Z��41�gq�I�e
��|sb���DL�ش���'oe-��?&�a= U�<����-���w�L1"�q��M(�l^x���DHOnt8
�z��a?��ѫ�����G灞��,����i�)�J0)oa*�EQal�Ij�ʟ��+�B�ެt(t*��KN�+�N
�q��5]��]�`���Y��`r7j!Hv�b�EH=�u�1�������j��vx�i}:�[�QGƢ�Ԯ��_��m������@lQ��Кr����Gh�,�z%T�u���0؏X�
�G\)j�o��q�� )�,Q����oA�ּ`Ŧh} #�v�$�n�L[��ЙCQy/M��
�MP��;^h뷞�#T�U�Q5e1ns>O�DV	�����]����CG[t��Iq!�Ű�L���!���1�"IU��9�xU�Y��-�|���2�1'��p���K�[r H<���K���ψM$��w�]���EM���]JU���ݢ�?��!�"m