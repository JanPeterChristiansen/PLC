XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����w⍡����,3��9j�y��Y��2?�����w*'�|�ݕД?���p��>&Sin�α����f��o���dr��B�
� [|�n���B��Q��4H��;O�=q/-3bQ8rS?ɶ8�ֲE�-�m�rs������W1βz.���G����l�@qOv�b�(=S7��-��hKKB��e� ����'�� ���[$[�wm���o�0KԜa�.L.˔("��d�w!�rT\�<��V�}��A&~�7���?!�� D�>#���p�LF�Ҕ-=Z*�
8̟y1���:�Jz?���7r�yM.";% #�s�����s���^K+�Zޡ�ܻI�bjE�w� ��y �kUy��������4右c�
�1��~P�gvw��:���ʬ��Y+.������7W�D��;�j��o�J��P�C-�ۗ�ۡ1R���bйB�i�KJN�Ϧ<�K��8��GF���c�B2(xL�RC̘ *Ӥ��,
j�>f�;���:Ҳo"A�y.!�����[����t�D�c׃�_�ķS����i�8p��ŏI�ol�����E A)��.�!�؉�T�c"t�pPNt|�h�7*ٕ��h��8�}#��}�W���+#~��"<�֟���Ì���~r��1Dï�^�ߤ���sؼ�Sb�q;������_TZvy�4�i6z�� ���p�P�5d��!YJS~��9��;H�c�:���?A�R�Φ��j���~�ATz���is��N2XlxVHYEB    56d2    12a0 �xd�����ټ⠅s@D/]��:�9;fy��4�����_�kh	��8�%�M�����eQ�x�]�8���I�Uckv	
�44���vB�w`eN7�����@M	d3�XSٗ �4���y0Bݰ��R��޽��u��Ҧ��J)��.��o�;@�Z��� ���J�����fO�`��E�I��g�DX�H�J�W^{[�?4�!!�c�4����RWHi���"��:��#Ϗ"\�/t�r���YQ�	��Z�KDb8�W���Zcr\��q6
H<sr�y���!m-��\�x�7�瑖��	�v�C~_�\IJؕ)]�aD��j� (��L�]K���p�;���L�����ۘ���?���6�MTKtp�46":!��_��8ne��W�u�k�'�n���~6�-������F�G+ ���soӵ��0~m2}z�ň���"�Y Q�;���v����F�'�D�+ ,�9 �I`��qH��}�X?LC��8I_�Îm��?
�Ep�V���GDmh�F΋cn�F�1�����7t���%�,�E�`/�@̥mù��Xyr����~� f�^-��a�>A��]f:1�LgA�kN�/
������Wj�� k�;T1��Y�D{$QQ�^��)�=_�̧���6���٬D$�*y�+���$?���Е�!�8��$G�A8��J�A+�O�X�	nd��	5�eb�q��4�����)E!@0n����{�Thʆw�D;p�2�P��!lfK�>�wp��:�A�������'ߩrq�.�)
������o�w��k�w�\�a�Wb࿠zL�~��R�>���4���!�z�S�������F�����Ekg-#�[t��j]8u�VE$:����7ph�m��Y���i�s�\�?w��1���+M���F��9~";&���3�5\�5���~�C�����E�:��q鯼��u��������q#�^�����E�3
�q���Ju��v�\�%�3�'<�*E'5�'ث����"e�I�/Mv%���1c�3��=�Ģt�	�L�ղ3��,+�t���Ci%G�DSy���8����� �v���|qC�����5��.�*��{&Oi�_�+J9��m�M�N]{���p̰9-A9��E���ܪ/�]ݍ�&��C� i?���,L�V{��k��R~�aZ,���䋃'0��Lp�C�1uku��m
��F��d}'�O�����1P?�mCl�u�;8�,���x�R�-_�=��r�l�<2����f�
��]&���A��wi�l�s�[�v��Yp��F�b鸱xo��?�����{�}Q~��'��O�bH����{L*?0��k�i�]%2�"[���#a��T�˱��>�k��=�Srˣ��ՁiA�sLU�D������%�:�Ow	Bw�3g�tu<(Q��X�q��d捍���J�^K�~{nK}w�(�VӪAٔ�W?3���J�Vԕ��9yOBg���g��lF����r
ϴ3�T��DN���x���r���л��������ҧ��=(ã[R����l^ja�\7�)O::f:��s�$-��i��T<�/�������90Xم�����hu�X�Y�q��f�E���N|�R����^{*6vݕ�Z�ËjD+�.Xj��p�E�Fu,��Ըr��
��K�R��ݛ�X	[O��p&6��}	@�Sg�����R��J��vϏ�p�T�ѳJbN���,�Pn��1���*��n#�N��jm�R�L,K�Z�c8�j���5��Bt�'�5����U�]p+�� �XU>�����N��KˮQ�1�ϽZ��އC�(y��Rn�a&�1kC��! �{س�.n����w��	�nS~{ 9N��U|�n����ɹ�`��c�ѠY>	o��8�y{��[a��K�a����Qo�����u[��x���l� �U�9vpU��Q��8�Dm�Y:WI��(�㾕�#</������gL��W��Up���L�#��)�<��+�[a�����WԔ9`�w$ۺ����I�����6�+�]܂Gs����P�F%3��Tp'��?�-�,�z�xr̆]E��y�~���L{�2�ӌ��F<�t������Z8=�U��k�i[�I������[
	���Ǧ<�5��X�Ma>,݉�C�9�jo�����!y����ƍYo�M��}(���V�xIn<�����qxo���GU�tn�g� �zi�\�Uj���!���nR.K�yx(�{���x�SpT&�ÜݥI~=���qaF���Z}y<o��\�q�z$��\��xn�з���S/w���j��x���'��l(�O W���Em,`&���0;<���%k{V��r��bXs�XPFm�Ax(�w:�<'��:��Kd�6�"8�8���m�[K���5�׈yl�XJ�c�����pt`%���>ۜ)���JV���j8�������d�xb1�-s�[�R��h��d�O�[A�Έ�.N����|	xV�v��T�4!O����T}[����y��s��q1�0
6���������b�������e�.^�^`s���~@���������)vvϚ�B ?��$�8*�FzO�>�� D�LHP��8�D� t���ٿe>vo�2�O��
\i�@ً�������d�E�Os����n�G���	��&��������sоHj_�*wUYg6��.�q�]k�[q�t�� Jl,�낪�4�+`��(�E�{�PT��0�O�T`����� Z���vA'�3~� �j�YY2�;��^�De�L�{��w�� Y�C�w�amP_�dX&!�
%\��e�fTņM!$�@+���Na_�s�.�Ӈ��X\~ixwYQ���W����w���}��xo �d֟$����[;�g���ж�Nت�pm��uqD9��-�uR%�:� Ş�Л[<x���@�G��!��x�|��\����t>X���Jc,6H��iQ�0�^�;:���$9��"�"I��g��XB�m[<'�O�
�-���?�y�kqq�$6�05��7FM����##�]C��
�fl�2�����,r�z�FVtN�̘��|�V��s%�@���W���޽$���k,�H��8�EK������f���K���)�d�eO�a:�G8�����J�~n{��[��!PHo.���R��W5��,�Xy��v�����?UB�
l�<ݼ�"�[ҕ�>�c��z�뉆
�|�q���\�޿�/��"V�.��q�?jNZCY���+�!SH�Ar��!��d@[4~��~m��"�!�\�/�E�������-2��$84MV�6�ޔ�d�*���j�vht�U<	�H�ٸ��X���C�l�8������\������T�ʗ�\Q��d>oDŽu�v-B�6>_�E5H���С�Z�g�dJ�H${�J���iι,���@��]G�h��G,�I�ϵ^� ��\oݾ��;.�뎊_|�����TMW��p K���|Fm���.*w@V�s)����w��O�SϾ���:b�H�݅}��^�kG>�"F_��'9���8���3UN�5�|��%[����s���CV�h�����~���߿��Eg�/�l��Nj'O�$����inm�p��v戫�*ϸ�⺌L7��1ݒ�L����zS���W>wx�B�5[�ܖu�LYqq�'���-�v�&�0٠��n�)h'΄q/��pϞU�)@�G$�l�[Sc�n:cƛ���S�A�v���L����,�����3�{�t��`5��>*q8@����![��4���P��H�ū��W����T���M"@8*�עIb������l?��^u:^rl��w@-�
���G�r!���8�A�#vY��=�|YmV�)��^�����6���a���|�ݵ��*���X�3-F"����}�N�?�4�G}�@뤣23�}�+^��a�T��HC�U��0#w�d$"�h�@|�E����2��=1j#}�SRV{9I��0L�o��"HQ��;�d�� ����&$��v�q=M)<к�A���[V?u���J�k6��2H�s��'3Eg�Z��@fa��G�� �Y	W��-�5��]�q�Ҁ�=ٕ/'.�����p�bj��`�Y����:�ZQJ��q���#�J�ϙ�3��gyC/���l/�xc���+��Ⱥ�ߒc���-�h���O$��7%���4�U*6�>�/�,��<���[�}�.��Q}c�r	�):��q0	V@�е���?F,�*R}��}��8r���ҙ#O��?��,u#��C['d#\��/� ͌u�r�4^Ө�o��am%.����N���d�d>�p����)��/U�����������uwQJ	X�V���0��|�ˑ�5̥{��l�s���D���)��'�Z��מl�v	S���MU��/-�Q7�/���In+����}�EA��:��ri�˝��ֽ��a���� �`� d�}s��5��IB��+��.�6E�k$�3!O�9\rȒ�f����5{��T���ܕ�@�'ap%�f̦h'񇼪�X]�