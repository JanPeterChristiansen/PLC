XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����A�|�=}�\����/$��3��I�����ş��|��YS�1u���^�o����)<����;Xխ�*�a��� n볒��rxSF=��_O$&�ղ���اvV�f;bR��0B7YҿO�*���5Y3~��**d�������E�±b���pD~�9�VQ�BZd9��,gMG^��j��VU2�;��'�o��݃��Q����,�GN�
z@�{J���(��Z#����C��pTd��llR �;�g��� ����P�,lR����X��&�����`�������X������ZC� ����4`���g(?�P�~t�h.��p���2I��!Wֿ=�ev�)$�
m��c���!F���|@zM����2ڎ��G�PX�cO��:(tp���8���|"� ��W�S��J:��KY#����_J_9�p�!8��D��;�pld!�u?h�a���8�x&�,�p,Q�)@f9����.��8����[�q6�A�ͅ�c�Y �coIr�x˭k�5�Й��R�(���I`��ʗ�[�+j⮎���V��X��iXSX��B_+¬M�BT�W��p#P9�2d��r"�!<6U�w�r�'t����"����*�,�D��6QQ�Q�f�,�A�����oC���"�׍��{ѣ[q�?;���66ӂߡ�ρJrMM� ���hҵ�������㴂�����?�����Ws��=�N%l���q-��b������w��󗅲M�@XlxVHYEB    fa00    1ca0'����qG�����#�۷|���Lim�M�����Vlu��]�C$$4�_�¸��L�֦�ה���[m�J�o�f�m㬞�DE;�DhG�~�' :kiȤ��9�&(���6�KYZ�J�]�8!�5�ȸCtLR�/s7�1�Vb¡Ę	/�S���'��)Ǉ"m�����w"���_jkO�iW���1�G��H�bC,�J��Fe�`ߏ:O�(���R��/�fM�J�둻<�~Y��.~���=�{7��W�1��Wr]ËE����Mqאב�Go�
<"�
F�g�b_�_���k�i�$c8�E�������������z
��P k�~�,/��v���gᦜ,�xf�\+P7��+:�ɏ��5���d�8mc:sL�hPډ�T.g1̟��`<ޠ��u��������qs7ҥ����qq�š��O)��lYX$����;�E$�u�F�e ���� ��Lyz��D���"�O�U�2ą�mR��5k�4�n�&�х��̒���n�	�k�������C������C��_�,�m�lVD̒\CH+ª�y �K������Ӿ��qt��3��=\q ��xʃ�C0�y]Џ�r�w#H�_4��'�������#�P���CD���T`�2�r���[�%s�.R��O,�w�U��a��1(Y��L��Rw�Ud=�r�'�8F�q¢��@��n�T�+��S���0ni�����:�#B2�PD���O~�-��y���⁜c��^Ф�3�&�z^}���ѫhj��.���M�s$8�N�⠼��HaR�N�PblJ�S2�)NV�u�\�|~Z�yC�xW.�r%��M�v��4�ųW������Bj�Ƶɑ�T�x�4V���J�榄�jFaܚ[���nYd�����Xlu���UA�%�j|��a
�]���UAp1�>ʶ�BPu��\����/�
�_��O�a#��B��!|��,k�9�|p7A�k<���FT�5̏&dL8\�eKWX�bn �]~���{�\�x�ٜ��A��mG���r!���)��D��<u�E���}EV6\��.��#�1��Cܣq��q�q�8�
 }lgeu�I�E�c�AI��ȱ�mВ��$颩�����m�	�C��f>��ߋ�T�z{G�ud��a�ɀ�5��Ri�Or�@r�4�wU�U�y�.Т�u!9�B�	#�H]3����l�'XŴe\�Tʨ��R<�RTv?d��ZU�x��,#V���%�z�jf(��'R�#�'=թ=&K�q��r������x�m���/�g��҅�@�[�r�!Vp�sA�-�vŶ|@���B��#�Tl��U}W�d��R�A�o�WK��[���7$����oMJ��T�Q�6yK� $AI�K����N��M����<�EI�]����/���֍��M�G��=m֪}ݻd |��A�"btQ��_��Q�:�
�})&z�-�9��%ř�2߅�g�õ�s�� `�]PdF��D��bxAt�l�o��x�I��H�#���߳j>DpӇ��2����%cxE�Q��|X����k�P1\dJ�ǥF=Sق�|+r(ւ�M�ܼߤHW���C��2�>��R�L1��4��p���)Z��?@�$�V�ڑS�.��#��T��ʐ�<��kqhh��˨����H�f�$Ũ$v0k&����ȱ��l�����0�/]&:e�������Y�Q��NW/��Ò���3c(�Ds��٘T�L��� �/Es��;�[͚�B&>��yd����y����$~V�;�3�S�j�ΪB���m����¦� r�џ�t"����l09��N�y�cF�t����]�<��Ae�,ܱ�k��/6�)5
�9Ӄ��P�o�x�L�4;=���9���e���El��Q^e3@��25��)B0�Q�]d�Y��:hF9ԈB��b������שbM ��F�$��~�����:ֆ��
V�5J̔^v��W !V�!��L&��G��/
���v��:��qX�Q!#�S�з��x?3ȫ���Kы�z=��/����m%������n�J�����kZ�F3�æ�(,�R��9d�8�h�u�w��L���*��'F��k��0_z1��*&$I�5��g��0%u
�PZ��$ڋ_������/�<FTF�ŕ���S���u~O�X����#��W �b�%�Y��������*-` �Ҭ�눨R(��ڳ+D�U\�Mu
.R�^�QW���["��S���	��Z;b��� ���@i+|Z�yD�%5A��|�z뇚<�9��2봃O��s�/�;�_�3q�pu�5'G�B����CI��}� d�-c*]�>����k�(���X�p�V'Ej����KF+m�ԀӠ!� ��]�)�ȿh��_��ޢr���kc�V����f��,��ː����G��n��v�<\3ye��E.�K)���3Po���'1x���/�ɰ��݇��26�]�'��1'�GB��;h�e�A>��B��u��J�ja�E���(�>k�U���f=w�p)cMh�1!f�����I_�n�z�'���*���D�6�Hh�9��VF�(�X��Lz��l�0-��C5�e�Ld�]^�á-Vt-I_�U��g�[��,�U�_^$��c/��ѿ�&J-�&��O��E�QD2�g$-�rİ�pO.�#2��HС��zq!L�1��9צUh�7B���~�օ���9u:D�����7}Q��I�Qj�=��q}��<y(��㲜f8wpM�f��/��\{�S�R���K|G�-'�+�s%F��w\a �5��mN`IK�L+���)J�J��T4f���$�������#�Cx���8���BFʒӹԻÛKG�$f����8ɍ�|ЗWu�OV{H[A���aX�(���N���
]�ωE��S�����E�T��l��Y�B�����\�?LI���t�@+��q�pLL�d�b�,M�y���\���HZ��Ph��W�^����z�5YKp��I�c�A��dk�������Į��E��v$�%�l���l�W3��!�z�
�3q�JN�/r�k�p~H���-Gɉ�F����od�T����~	�O'�þ��!NL)q�*V��Jr�ȥ�T�gdXF��� ����NH���vk;?�|SVC1G>����<2䮵���U@1Ot��p�����|w ש!�Y)�D�[��� s�)[,�\��K��Ym�SR�.Y}w���k�1�����FGrr�I�Fc�9iXT+����?Z��/����2��*�"EqŖq���A�-� U��w0�~�*p���a͟t$[6��{#{ëLrV��8��1JƔ��2�E�)3�9n7�W��(8�����#e��B!�͚HT�بRkA�NA>'�����ڼ�<���cm�i'#Ĭ�%ĨI�ѡ��L�O�IE�Uw�d�� ǐ���W��dҚ�7zuƺ��J��ׅw�g�3�@ͼ��>y�DH��E��")�O6F��X��9�a���Z�N� BC�>Z0e����4��3)׋YRS,�Zv-�H��n�ֶ<����
�3��6x����Q���rOo!Wܑq���$�"u���<n�F�}��[�G5��s.EĎ�)?2��	s���P����D�⎁K���,nĹz.�~�d1�I�SC�5����]L~+�� �Յ�F@B���B��`����|fI��J�A����C�r/���_���c�͊�.��qF��t�ѹ�J�<�aDf�*��Y��`B��	�H�/�ׯ:�8���a L��|�CMu�V���nf�wz���/w�#Z�٪x��|s��S���܍����'v��l)�y|����a懗�3�(�ê��q��kI�X�ߜ�Iw��3���?>��^�~�LH�G�]�o�	��q��ͭƂ<�SF�>���4�[uDrbSxy�ϥ�(7]9a 嬏v��뻭f�=9Cö�[wމgw U����s��0�������7�e�q\��E�!?��*�7�@�7��_wŰ��G0
K��%��ʋ���J��t �֋�O�_��nm��)�	��F�ܭ<�s�-0K>�a/��܆��@�h-]��P�o,h���"o�P���[�ti��Y��� ��޶͝Y7��X)����z�I��2��Z�-ߵ'h�H3�A��;e���T�&~����/��J�O9?|mn�O���Q���>��#/�4�ۺ��3���]UF)�m�j�1x��Ҟ�z��I�=��zZG�T�T}r��|��b��sЙ5�$@%���`td?n���v�k��D�N:O� c���X��ܣ�Jx��VQ୒����\����I�Q��ޒ�H��>��5�}��WD'/�s��d��rܳ�#ݰ���&���e5�õ��r����� Q�q��CCqc�Ŕ�P�����AB*�?7���]G��pf�?�a����b�j_iI���4��%pT�P ��������9��1=,� ��(�;�Ԩm��R��1�@���^�1��rcn��4�=#�B��B-��u孽�<��~%@n�i�>%	n5��_�8�̱�t$��v�[��UhZZ��<��Cf�sn5��Q�IA@�3=�P)I��������;�{�Z�ɝ����t��0��(��4�n�J&w[~���&��-m��O{%ekiƩ2�/AQ:��!����2��n>�g�sX���*x�Nj� \Kto3���Dl��7`����A�镋Xݛ B*��ڢ��Е�icmN�b��n�{}��<���F�wD����ʟ ]S�ж����e��mʹ+�8e�ҋ0ӐwtF1�����F�٢]+�T%����+�y�&aF�5�s�6�i~�F�0)N������C�>�1$��J9)�
h���:Ŋ��ڭ�$�'�%c�#i�'���(�@�5�`|�*Y�k��)Xon̸�R���p ^�r�rK�^��;��@��&�$��:Ɂ�� ���5�PýI�E������3w��}Y[/:>�It+��I[/�����4����P~�-���C?�-�z`�M ;O�J.ɹ$R�lww}w|����Z��#��ἈY��4}F��)	�	>)�(����0 �� �QP����0����ֽ�9ف��
�߅����f8��#/~���?��4�&�Ӧo�Yl1�+�����8TJ�	��Dc�7�ͯ˫��Z|Bќ�����L���ڛ�!f�j���sjg%�����Ѫt�d�2޷������a4��i`��͏(e�bŤ��Ml��z������ ĖVtߦ{ 1��!@�!b�>�ɞKѯ3(K�栊�i��,kn�eN��Ro�^UL:����Uy�L���p�3�̳Y��=��'����:Œ��$$�m���?]�T�x6�6�f	�/��(n�M�F���d�L�P��^�t�0�������0㱥8��I=�L>����Y�x8�����(S�8	�0)c�dzJ$�uC�Tt��E1`Ju�߮�PP~	n��vaޜ9;p��{�!�����#�R '�CbE4�E���η�+HC�W��(qû�S���FT�4�Sc�Jv�7D�$��RH�$2_W)M��.�/�W�d�f��'��}�"hL@�t�굖ar����i���}�GI�?u��8�hj�����},�}���=�aIR� ���E��~�����ȳAe����s ��~��b'��9t��W�5G�A�Q�9[mgI:�*�S9j:{���q�lOG3Z1�~���R��ꮶ��b�1zKeٜ�� ���Jf.p�+s%��F�I'R�A��Aj�'�uZw�he��Z	\�{7;��'Jn�z��xЋ���� �9��P��\�E0T�H?]��e�랖;��u�j�~��h�.�W��d1A��� �D�?N@tq&[ciS/}r��|���E��zWZ((�����vG���W��2W;�ϙ��)^HK����syX�܋�BS���.�k�&>����P���W�.Y��sfu�8�s��2�j�/�Ws��J��U��� �bj��I�R�e����O�*]
E+ਹOS?�*�VSL����!�M~�h���(��ߩ�[Y��)wέbC�G+=>Q����r��^b�Ī�5�w�����/fq`��a]�d��94�ڤ	����P���sn����F�$ 2���
+T��	�hG$�רu^�B��x�<�y�;�P��Iۨ��se�"s��u�꥚�E�K�`|�y.!`]�Yi����M���<<���dv�@N�=�9P@m��_MT��h8�Ψ�w�<!��8�&�i��O� �J���9�Gڧ���o@fkD�0�,�!'��{���,G�q\F(�y���#���n��f�x:��^��.!��Ų&Hߜ��輪�z#TN�Īw��VI��ʞ����Ӗp�SB����6��+���#У�bk/E����W�l�S��U>����� ƸBh����y䣗b���t!P1�V��X���kW };�G.����"������cLM���hnC����l:��M I·ݲb�I�cB��&����=��̎5�BD'X��B��#���Y��c��?���Y=���Y�[��%e���wZ����HJ��\o�B4�L�T�T�nrKA�j�=oalQ�~���ȱu�"v{��\J?�\c�}�r�\�_�j�울�!�1i2-��P����ӗ~ �&G,-��5[�%�_aO�y � HΈD�]������T��R����P��^���=�����^ �7���S��g�,6f�VJY�� P�����V|}X�z���_M���㾧�� ��h	.]8uJ��,�)���À�KD� ��}�I<�(�v���\z��L+-�_�P���q Er��q���a<2��[�.;�?��JQ�i���,C�)W-p���5@�S�,`�8�F�s��o���Ɨ]D�.��l�]�f��z�])�56���ȳ�dC��jn��q���G�v6���dR��F��~R��7J�}m\W�1L7Oq4P��$��{�7$J�&�97�7[��ݺ����b�dL8X�F\AHI����Mл��[N=��?U�$;�3�z6�ST�i�fM�T%]�"/�.�>]n�`@���w�VO�Q�ȥ��M�cXlxVHYEB    fa00     cf0��GK���8����uc�ʌ�U4�}Φ�$���M|�OŢ�2p��:�)�����X�?�&���$��*N��X�Ԩd��I�L���� �>zL��������w 
pVc��S]h�%��q��[1i)��?��%�N`�:�a.���Bn*�9�0n�x�P-��"n\v6�'�����0����AI�O�a��:}R��m͘�s��ܧO؅P3*K��&=�^d���C�߿@�z�@�f�����rAW�QZ*��$�wu��va�h��(�:�+����n�SD��4�d)�w�0�Yٽb���\>�Z�8�Sh�s��x�<ƛ�!�j,�/����	9���i���mJ��
�bz˽t#Dߤt$�x�8�S_E�li�	��St"#̕7���J�9�	y��>��1�T&&@M�	j=A���l3�qB�S�J����"��CR���������E��}Ⱦt�e�g
-���mlͧJН~@^Y%�ړwF0|�K�_�:�/	َ�k��cu	A/�!4�l �k�3K����y �m
��^�y�W��O�?Ƽ5[��>��2�\�>�l�n��{5; VBz3ʕ�v��)�%rN��5�%����#�o�v�0�Qz�7��_B�5�	�����1T��F�̓c��Ucq�[�OD�n�0Y���+=�H5��f�|�O��!��� ��7n���sQ�.N�w��#�~{��6y"��F{n-(6�r�>�4�����L��1����{E�p�0�\���v��2��	>< ~�H闪u�tA�©
���ojS0�m�#�#(hC�p��
�;�װu����B�*�l���d7����<7��( '7�?��B�î�d
$�y����v�p���S�`��F݋N��� ö�7��F	�����~<F9:�T�GM�xw��!����ڤ�W}��]E�2�|��ٵ��fi �`|���/1uө�gzzq�"���T����>́1�S�߄lՃ+J��P"x�
�"��2�����] 2_`�uW����*!��w>H*��
ڽx{�p�atFv��J�~����&p�P�,�g����Y@�ܸ�Qd�uǤ�����	�wҹ��	+|z�R���	�r���*��cdM6��b�m{��걒D\.$ ���EP�@�����q�<H�{V�5S=x�Y��Xa=S���5J��K�@��KꇁL�@6c����3Kg&E׃���/��a�jWK�:���NO
Q���sߖ���VUd�������4zQ��p����w�[���ԕv%x2뻋�w�#�~>�H�G~��(91�gǉ;�d��o��_��fnB�D�����0��<�^�&b(l4tv�X�uz�3���:�!BP����8~���R�<-���Nkd�w��ba!�>`����O�����`��A�YAn��X5������ x"��u�%�������t`��
-O>n��-�l/�c�|�-A�Cd�>�wLҬ]�Vo/,|'���\b�+:Io~g��'SM.��S��iVF�ܰ�~���D(ZC�f5e���M�3�w�B�i��,��^��i�! R#��^��U���P,D�%�%n���,;�{�5����ڹ���Q܉�ø�F���y��H�R��N̛&.^[dvi�{���46~1���tD���6_�H %]s��z�,�l��̔zñE5����{N�u�`��[�E�p(V����.�wM�6�ݵM/�H��#R�2��J ͛T15�ݽ��U��h����~D\���wo ћ^ҠN��&<:�S���zw�?�9G'�����|�����Ե��`�j��~�*ȘI����R��#�)����xZ��9D��T�`�Ex����{��_�Tx���*8I��_��D��E ���1����n�]bOL+��F��q�k����tV�K��±X�]�Y͍�J��/�ޱ���J��Ba��Mc�^j��*.�At�;�= ���ńN��g�s��FIi�M��L���t]1���$Y�=�o�A�;��(�%Inx�t�	�*h�qw;E���ѫ}/������7�����z�V� �Yџ�]�[ߵ{{�����_���=����-؍����KV�/�i���X>��R�UА�úe^����^Z�>n���2�����(��}F�į�	�w����S��}�+L{4n��s��w@��$����2��c��k�)��X �-��Ih��%���ܪ�P}Й몄V}�k�ؽW!/hwabn����W����G	��nU4B�a���p��肣U��mv:!�xЏ[�=d�jz]A��=ӵ,G��?�����W>����k7���.M���I|d���AAK|h�[�vM�'#��ms���)>.2�k�R��E�E#�w�����8���F?����]����H>Ѯ��Fu���9 $�r�p_,�`\0�d��_Gqu�
��ǌ}�u/D���I���b]�<�KB^^HD�P��J��.-[�]�L���X�1�4�u�n1F�>ԽS2��G$s���l� ǉ�j���f6����W�˴�PU6���+qU��ˊ������۔��n�G}�a���� �iD���(�E�Xga	2�V�Y���=O
L2�İ�O�|.�c���Z�tm��L\�'6� V^b���k��et����á�pѠp�W���ϞHu�Ћ��xUuU��7\��識�I![:�+�P�n[+轅)�K�^G
Щ�?���_Br�r�
�U�:Pl��;� �Ww�F��Wv�oˋ�C���P�}dz3����eĭ&$n$�
��a����T���7�+P�m�G�Ku�T���?��`�[�5��$�Yϙ>�����fK�ҼU'L�+�g��byT`kX����&�E��	�(�
c�3�R���W� ?]����ł��1��@��	��:�	�<��y��|k^�L^�;r�o�;���}s���
]��̶>�e$I"	1�o�[.�U�H����ހ���j��Q��d
q[p�R�<�]˘��%<#��#�g��D�֓)S�W͏�������$^Ni��!빟Q�0�셒A$���^mw���T��!I���S��=*�����,qXc�o���T�����mrɝ�n���k���b��!Hu�V���E��/7edkwв]���S!��_'��L�y��Wz��M����Ә��ƽa[�:z��T�`��V?���XlxVHYEB    3981     4d0@QR�.�'��$�� ��ڍ���@@x� {:�������� 1��r������yt; !��C7����y�lJzåx�ߥNr�S��W�@������q9�1�^��&�I�໏䡸f�84�mj��ƈt�4R���Yx��L*���v����Ǌ�����D'���[ڙ`Jܠ�W6�#���YD1��Sp�J`T��WL�k�/�~�<��Ѣ&��7�0h��{>3���� ��m��Ѫ �VM���r��}����mpKceVb `�Br�Eh��O�}Pә��,��z�DP�7��&u�H����4bQ��l\ys�"�Pu�[pC!{���c���l�f]����?��TH�?���w�1v�;����.a�/E����5�ᵚ��<�!r��x͡1�ֶ���p���C<M�/B�~�� ��YE�
�:}��Gi�~!�`z��M㷯�%� ��xN�GIN�7�f��D�@��jC*�J��{�Bz��v�n�M��]����G�o}1��ڝ�t�;V}���|-^�됑sb h�"�fz��Ӡ1�Ēx,��S�����t�`���=�����F>�pLJ���Ӈ�T�2ɳ�-�=F*6���8}l����\��9���%�7���c*V(N[F���A� �E��n�Y�C5���el�?��Pi��h��x�v�bV���O�u����o"bL���iemXe�) �����n�Ƨw6��m��fT(e�a���QP�������j�xQ�Gb�.bC3�"O�X0�7�P����
�XP�dߠ	�f.��dC"�ԧ8�����D���T�+F����(����u�X�i�lV�.҂N�N
p"�F/����iΖW0��ڑ ���0M#k��:���A���p��Nl���3b+��k�%͵�ȭ$���T�ypN4����CN��d�M����̯�U��v{�k���ɉ��� �����e�~%��lM=����4�o%���r5�p�U��d��BR�Nܧ,O��R,������C21R@��i)��+�s���#߈Q9��~J���
���kv>����Rs)�.��u�6�ɗ�'օ�܎�.�a�f0��l@�+-��s���������{�~;��\i�e�.��D����LL�����vd>a{ѱlD�����B�� 6��1
  ͗^��q���|A����!��