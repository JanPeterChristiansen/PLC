XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���/�y�kfIr�O	�I(n���ܦ���X�[y��U��	�Y� �S��g%��D$�Yޞ>�w��� ���>�p��W����-��:LN���������6��L>��~ ���rO�M��j-�0��{1�0v�N	�2Y�du�}�S��:�y����ɿ3YF�g��Q�e�[�MJ�k��)s�ض��Y$���]`B�r>l'o��P��4PT彯-7����U�-]'&~I'|�&���|�{5KBɦS�"�tR��_Ut����甇��/��R\o��#��ZI~�~������Y������>�\���\]��~n��db�s�6��#���-�
T�ox��[����wd�S��n��Y_��x�K1�<Z88�	;�/����8b��+���۳3�
�(��b}
���a�ɿ+YC��bU�C)R�Ω�7����떼�n�c��+��z5R�'�2�K�%�Ҭ�^(��i�{��t�����'Lm����Y!�[N-�-��ӳՀa�����CFz���m]az����"����k��A���R\��c"�H����S�f��6���3QT(Y�5 Y3gO�K��l�y�z.m`��S��R�7`~�MSl�ωz<�$
~��z���^�M �hw���r���/9	�AZť� }=\%��:923��X�nI}�Ch+p �Sϱ �!�)�g`Hӊ��z�t��H���Z��z�ַPB���[���d��V���~��@+/��lXlxVHYEB    fa00    1fd0T�w;��.4��e`��	�g�;Կ���o�\�_�B;��.���fXED�N��*Oň؅��W������w/�D��e:��E����+f�}i1��q�5j�J�S#*���6��iθ�Š�B	�3,6��o^������ Oy	��9@A(Y�w�{��'��qh�a&0gD����WT_p����p�L�(;���d?kJ!����O��#)n��h�:�ϴ/?�Á��z��H���}�X�����^haQ�]��1�SYkS��*���ʺP��;b����+,O9��'��N����vE�:}E\����zs�p�iC��}��>ۘ0ɯ"7ͽ�2�NWJ������kD�Zi�_{ZA>�����p�\�}�b$�:���l�2���s/��q����d΃���f޹;�ԛ3���CQ�V)7e���a7��7�zzb�]N-p.���v1ch+��#���x7�dpqN�'d���%�&k��j�EFK��kU���s;���bCр�Ȳ����L��'�Y�C�:aroBo�,.~dkU )�jd=nd�}=Z[���3�3sT���Z%������Wa�@�Z-����-�	U(��S��CX�qPy��xv�������,+�O�;�ʏ�Փ?�m��#Y��b�G�C� sP����yZ,�ў)>�L�P��^�:��~�a�͚�Dp\�u֍�^�]����?Í>�q������)�m�.�;���J��a�Z��~8o'������ �>P}ʇ����B.�b0er�2{�t���ݞT���^�5��H	�¹���e<��>(LC�I���F�Y;x�������#�X��a�Ϋ��}��J����������L}9�uc�>�ؔ����ϴ��r�t�8���`z���iv��7��u���PȆY�p/� ��|�@�mc;)�i�o���W�ȗt��RH��7�7��i�	�ǟ�IN[,�ˈ�u��h���j�|��XvW���V��y��a4��w��k~Pc��_`3�Q�?d���"�: 9�@;� �R�!�Q��Zr�ā��C�a5R�U�����̈́�M�O6m��k��2�y>+��a�z�G�GD�s�+�aE���/I��W�*�f�QA<����Dwu�S���P��Q��~h'	�yBHc[����$H>f)Z�˵�2u��w�^��U��=����H���%�lb��	�����| ��F�:J�a҉a��@v#�%+�/��sk�u�:��s:c�S�	��6�}6�J�����Ͷ�p	��{���:��Kf�����l�m.���G���VR�j箸��y�=���9���"����Vu>3�$|�7\ʿ��O��z]�K�]�i.|t��@_nw�&(��H�&�|X9�����R	�RJ��M�uwh}�.������	셿.ZѳO3����{u�Gg�J9��ݘ'��v�*�z�U�����w)_�oA��L�Ё��ױ���6�x��HZ]N��z���1?���g�$kHDޝ�)�3�h� ��&���C�ъ�]ۼ��˭�wG}yZl�����ԫFͪ۲�s���%6dd��[�OK�|�!v7�H��q��K��'�F#)�L��"�N#6�/c!ĽY9�!A���|N ky��P�BOs�j�Ӑ3p�
�΍�!/�Dp9�q��;�@�m�.��jrS�?��[�D�&�U^���H�{q�t�x��\�{�7�4�FlqCf]B�\/h}ܙ 1)�r9���|�QA�B��W����5����>�xl�h313�*�u���W��3�TV&��{a���م[�$I��Oj��5�搼?
��s�+��e(��(�.M��X��%c�;W	"2
("q*{���rgs�M�j�W>Ri9�.C�mEg����e�"�O��c7Du208��ER=ìW�
"�Μ���ي��N�ĵA��\���ԩ��a���Ĩ�ݙ�@��'~M��h�E����C�2�����n�EOz�v��<P���4r�.�>O�e'�_��W�A����4���*=&���Ƞ7��+�,89G��CS��	�����^x��������R��=����/����$w4��^�E���^�{��?t��}�oꘘ	�K�zѼ���#�	ˉo�Z5�֌��Ų+����濟���~jN��*�oJ���u�>�w�'}���߈��nCp�� �㦼���,�&20v�!E��e�b�2
k;�|)�Ŋ����j�;��1�Ss�� ���`|E���8����FJh�hj�������:I�9��҉�i�K�C��(���M���ۆ\_��4f��y{�� ��b���4�Ъ��Òf��#�EߊEq�*�:�H��0�̀��0����v������#M�5&X�ϡNN'Fl7b�9M�r�#C��*J<9ɍ���̩9�zB�B�E��ӌ�E�H>�>�ϖ�^�MGW@�]A�TI�s���̋�?�"�!�V�ʌ��o	.�ֈ-�v<{�o��33�H}��N$�� �xL�U����݊�Fb�T~mɥ�dh%��O�5ˉ�wz��'Կ\�}�Vx��Iuy�<W���Q����1a��ݘ��睻�n��zٮ���e��%�eg<�|�L��bwH�	>T�|^���lu�`?�� G�q�d�p\~��?�L!�t�H	�c�w�G�/;-aU'K�=�w��_GxFh,��,cJ��=�XP��ː�b�����,֒�	�e��b�pr���W��+��)�%<l��.;�b��><�R��b��4�4�N:Y��|d�-�U�P�bδ��T�~!?�ݽB
����o�ܔ.��l*l��mR�N0�/�(Sb��F:[ j��{���[BV����"���ц
J���OYy!��I1N}�)C�'��^�F��:����F�)����vi;��|h��Bx��� 'e�]�8�e	� �P&G��U�~8!&sdL}���CjJdo�geAw2�d�T�+��c2,�R�ޔ��0͢LuEM*X��` �]i���c�Z�"丧4����N�)�v��wAy�'��OK���%2_)��s�W\ݬպ�ἰ�s�ۉf��{!�e�3y������*�>=\	MI�;��g!�B[�>%�	_2�Kǹ�m/�`uz@�

�����?��z�i+3&{��q���Z*��u��0C�r�׳���?� �,��;@���<�c�'T�zʥ{K�cfe3E{�rm� ��{[����ȿ��&V�]���#��Yl���dq-R�S�A��Iy&���:u��������}G`	�<�!� x�q_Θl��n���Mb�;	 ����y��|����Ye�lZٳťȄHzE����ws���@榵�߲��1��7�(�G3C8?��-c��\�dx�xM�8fO��?Jȕ2�h�DHOn������(N�^�-�c/���v8�t_�e��z���d��|�Řa�G�8B@(�~i�ώ˥Uw�A{�[vM�|�~F2�-M����jpӯ��҃��\���t�p��C��$D�3`�3Ϝh�g������A�d�W��)wT�}��A$$�Hd�S�O��Htz|�����{��B�+=jG\9�tAYlqn�/���i�[�N�(�PA��l��<�d�嗯���R,6�eyvβ���i$Ս�:Y/�mC/B�L];> D{
�8��;��?bd�FEq4k?�����W0B���u`�x�q���2l��s߼�An�}Rr��,�[t���UדG�����>%����8ש��>�`^f��ҫ�<�nQ�g����gT��D{`/��1����i���C]zc[&/^C��u�mZ�w��	�5�ҡW�C��C~���N�������3eڹam��l�V�����:�X(s�d��`W��6=�6LS���h~Q���(fk�������'��V����}���&6��qi�?:��z;Z���U�d8�?.������ ��#/�M�my�~�_�o#.��G��p��X�&��D�f\$! s��c��>+]"Z��8�������W,�	T�$���>�r픾�#NyF*��6�Ŗ@��I����Y���`3��%�l���T��Sb�Js;(�h��=�3���̮q�@�k|���ms������7?�O<~M��c��L�޶zm����Fc���cG�M�{���=���y6��d=���o�ZǀGc�@d��B �ji[{/�)���]i��
	wL(p�����CfD�[����h�Uލ!eŶ1(4���qvv��(Z 6�Ҋ{;d��ì�w��ŧ���1Fs����(�J㸗zV��>"	����XzL����������"<�6��~N�#Y�3�$�8o��$�RN��)}��H\�@��2�Y���΀�
��7m�P(�E;+<�h<E0���rt�����N.8H���V��aa�sJ�%�j�K(z��d�Jp.��Mxp��`sh f��TX��S+~~偂�%�B����3D��͞��<���o��܋���F^�`�Ѵ)kF����W�m O@�jxm�����$=��@S/\-g��]�V��. �W��F�(���f郝�w@�ʏ��֞��J�d���v�ࡴ<
��%��'׎�s�N_��,NJ�Ew��i,c �-W�FLQ�{iy'a:~Y&���y�\�J�C��e�Ӻh����3��,�6h�7�AY��H��$;=3C,	�]N�[r*|�Ե?���a�uml�W�3�2������2E���Fm��Z`���9�zdaw-�����h�>�K�O��{\(���/Q2���H������Xyfx������-V���N��	� ]T�-����)y���(��Ӑ�����5	�tLq�[�C=V���ǅ%�NG���i+� ��%x�IV�y�E����n9s�gd9�u��U?�
�)=�9���a#���B�0���8<&4��$<��sWkehu������%��a������� �(�Fd���#c܄ |:�?!�؃���w.�=m�}i���G?u
@�e�!�z�F�O��VJ]I*M��q����5��1�s��r��`ȋz�^+�#�g��ܙ��O����~m�MDJl����p�f����xҥ��d�&�\���F�X�,.���~�T62��]�Ţ�<W"8[�F�t�� ���\Bh㈚�m��' ���
<����Hw�z����1�Bd���)Uᨣ�IM�B[�Y� 	~g��#uIV���)fy5ew�"/�s�8[��ڙ�5Vʍ�5�7hV�q3Z��$OV��L�F��4(}�����ݐ�T�fE4�?)����P\�2/�Ax)lu�����XDs�J"��d<�o�Ѹ[��̜�4�ɭ���>9r(�T"�ĸJ�Q� ]��Y֮��!�� �[����a��}����y�)ͮe@�%�������@�"v�G��~}���ȧ��r��Y��Cpnnݑ�I���<��R�v0�շ/ �fpR�N��Pt����e�X ����^Y�w�؛lو�����=ƌ�K��B�� ����ִ�\���2O!����8�Ɣ�\}� e �أ�G� �������o��η׬�!�Q�%�}���.o�.g����k�g��̃�d���>^������qb��ߧ
��2L�I��2�\��Y(�T��M��dmd�	�#�qA*�ת���B̀(
���p����w�﫮V�E%M��:2׼k�0�zȉ�*bT[��K�!�*$(�F�2��xO�iZ�Z�Ĭ3g��d�#��n��]㇀�p��"%�j4ȏ aH�a���"�&wՅ�>�q`Ju4����\Y�ïk+��kR�{�5-�`������4@�Z~ܜ&}�SB:��r�_oO׉Sf���0&����!��Ф�{ ��D���L��XH��'J_̕%������9<���v�{��ufGϺR��M'�Ǫ��jyh�y!���t�[��Qg([A
X��0�>��w�
�'|C�[���h�<|-U.:��؝�"� ���ݦ�o1طvYn��_qR�Yc�qp����@�|�2�|N��=V��<^��^q_M|9�#�{*��xi��/��#�Q(;)���WHG��uc9(ւ�-eѫQ7�S�=e�ru�lN��U�e�3�]Ǭ��"ɽ;�b��i�&52��N���� I�)@���{t�6��&��>g�j��ytM�f�-��ÌE��#���*L�EOJ�W*�l�`�/o���8�G���=������;��헀r�ߦ�V��/|�u杘��f�:����|���/���A�F����uޯns�f�z�����Tp�`��E ݫ�`8����؊�T�zm��ӽ�Z�x�sOI�"�O�U�m���sc�Uy����AHݪ!���'I��NynG�O2��#)!�l=��<TP���V��ЭU~��-
j͗j& �t�+�� �73U�a��[��YGe��7�*�A(�e��(�SJ�F�UZ��j�Nk�A����4\ҷǑ� y)g԰���Ԅ>���18�p��TB��<�-�"�\���a%ز5T�]O1݊�7���b��E�e���#�hM'�x�t,�xZ~>Ġi%���`ʜC���^̒��L�0��mf4�W�O�w�vi\x�R�Á��]]�0e��x�f��/'���..���ߧ�Z�����Z�����,��$@;��	�<K�sU��i�JA�>��%{l�:9�`�}P$��3ۖDv�8sL�Fz����b|�3/�jj578�-��#��[;�Ō�w{)$CG�(Kf����I���Y
N:)F:8�k��{�c�őo�����6wC��(�Ԃ�����0�/v����^��$4"ab�Z;��L��N�{��[Ae�h��=�������\8�$W5rE������%����Ȏ�}#�W�>O��:tد&������Y~O�n�,�\�Ș�2v~�ےE�RQ�-$2z�����=L�Zv9(�	�����R��w��V�]p�ŏظ�V�(�A񩸥�߅����}O�;(.\��x�ɒ���@�3J!�*���,�sߕ����nk�c��!TPH� �)�׆BFm��DfFNt6��6���P-*�̋3�#�*B�5b�<S��K���W���Y��S�14�������) o�?$� ʰ�, 8(����k���Xh�D��z����0;n�b�/J�O����bs�
��E���*���FT������a����p����f�U��4(��bm2|eӦ 0�)X�1TȲ�A����6��o���_�<�:�:���z���+�Iq~�̕3�X7A���k� ��> D�`�wTvW�^���RP��p��+{�F�y�ćH1�Gc)����&�	Ř����rم-_����`8M�3�/�N���܈1�c��My��M�/��ȶB��wk-�'P�/g��˂;9R�/�(�h�1ץ��V3A�� �pl��L����*JM���k7-0F��[��~f��]2v浔)Z�te�wx�v�3,�K*fN!G�^V����SR��SI����-�B�x1Q�zI�����)�x�tf\e�y������x��9o�t���1.�y^aP�g��t�p�v�ׅ����˗�����X�7T��:0Tw_S^}�;�����+E�~N� a�Wא�O�<���g��-HT��<�%�u�ϳ/sb}�lF� 1���gGv��s ��k�U���b]���$I;�E�Gmo��������h���̳��$ �,~e��l@��*Mʿ�������X_dd�ٮ��D˄�Ioq<}�a3�����bU6�i��>T�&���lc1�pmKf�%4@B	�Ǳ�Q#w+�Z9�4�Ԃli}���� K���㲌
��G�&�\��t��.�.����\P�6(a��6 �I ^隲�t�ݟ�cP'#��簕AT9ϳ-�qj��I�9�XlxVHYEB    fa00    1340[b[$��h��F��7s�v7��������ޛ`��ϻeWa��;��M���p�<�s��ߙ����[��'c=�~�1�E��M��Ė����-L
ٙ\=ڨ
���d�_#�Ϩ����8�>;���BH@q������������>�8��Kܺ�����wY(Ԭ����]��ڗ<�*`b&�9�Sr��L�p�EϮ��=$�u���XymбLY��d�-�+�d��Nc5�t�n���}˳�JZ���do/-���к�W���	=�g
�S�Ȇ��P�;��.�<��Q^h�V�@��HiES�ƛ�X&���˕�x
e"A�d��pQ跣3 �v20����ɱ��q�s�}].^�_2�rVl�8`$D�H�µE�%�q�;�m�r�j�[7 Q�+�M���_�ft�^�B �Ķ1N�VҲ�ul1L���jA���G".��m�&n�>�n�\�O.&�ލ<^���.�0��So���%�9)��� !���_��A���z��8���t%�ZJ�a��t�Bo'W��>ɩ:MEJZ�U9�[�!��=� [x�����Y���Dp�k0���U-���j��� \�X)�4:�t+:W���T�]2p�RP��Dѳ=kS/�g@���e�B��2ԴK���|��a��ߺ�1��
�OcZ��H����6ǋ�hx9r#���?���q�Hq�?��أ���x�	� �U�8o-?�B��]n��ae�y����Gp�X���Xlt�rrVz�S9�N�9�'��f+�jIf�a��7�r�B��$l��KQ����[/1���ޖ��y7{�t��9�Q���b/ �t�XM*�J�e��N	2��]�Z(�o8���1[_xx9Ҫ���T�M����W}BC�\�Z��u�|�L�%3P�$���w��q(l:�	o��6�eF���R`���Mn]W	ID��EFm�_�� �!��wff/�k�It"z�l���y�IΔ?�*>����<8.L<�#�16<f�;��#�u�%j̃d1J�Ғ��9�B���¾�P4}0�vC'T�-�����Z�ř��mIb�8C �ь�H���"3��dP�`�q�H�M	ф%��a-����ܞ�Jn��S��Z�!3��c-���P�Y%@S�{~�&��R�;	�VG܇
B��qwR���*�b �G㒛�	�,$gs�W�o6�g���kT��O��B�����T��£2�F�� g��0�N%?"?�/�E�n��'���_s}�����)��ߓ�o�3���C�7���QC�B�~�p�!�o-y�e"]�����T���~�XM�U͚��o;��T$�G^vE
5��u1ɛ�E�y?QM�p�Ӎ{��sb�~��Jɜ$�DU�p�B��/b�m���5�Z��ٻXc��\sN��f�u/w9�+��6��m>�w'�긇&�EK4��JM����<���0i���6�/
�K�uk�QW+�.}0�ӥr����NѪ3k�6�����S��\h�(�&��*'(Q�L�J� �n :=�^��M��m�n|G�pۊ{~� �iof��֛E�C1�
WN#�W��B[�"s#܂v��CY�֗zp \��hƁ��ř�TĐ,~��[������Н�fSW�"^�s͊�ߡ��̵��x}����|Y���{�fޮ�G�HQ#��p�\T��%p����2�_',�g1��ʥ��/��<XA�IMdh�n�?�Z�M�N��=qV�}��˒���.3#�#5�{��(��>�h;9��Sy��>� ��G�i�oO��po����ԑ0�pL���R�;�a�hwя�@؍'��ڹqv$*���L+L�ٛ���w��8��c�!�7���Ǌ����	�Um���1n>P���J�#\�����uQ0�P$�� 3X��Z��9��N��$8���d�ؠ�(�ʡ�@�Ǳ����.����'��ʂ�2)�LM��8~ C�PXbw�':l6��#�z�-��)��p�j��_n���H0�*�$����p6���E��P��+�7y��/�7�����a�*w��ݓ�Z;�ka����S{��24���z���yD��fDk@H��˟V����ɩ����jAP��`����P���!1�1B�5�A/X�q�
�����`�ZjCO�)���p��$��,ݏ)]��J���X������ZW=�m�bfO���v�!����e3�`#�i58�92ƪ�ĩ�k���ZK�PEB?t� _�Dw���p8�C�"~���Xxʆ3�·䑖Wv�T���	�����ⶒ�"��]���>�۬��L3�3�kU�_�0�L{]4s�Ѫ�+Һʲ��c/�A�7��H�4 j/��v��"]�o>�&��#}��w�_V{vL��q�Ϋ�@�`��ԩ����[�nͧ`�9>�ej��3�@�L���ړ�ͫ�@b�J�>���������V�ݵA�9[LmU:W ��f1��8��4�;܄��p}�3�!{D_l�sa	N��u|���e$^NY����Ō�CK���_j�s߅��ZP�=���Q��c}�n^e$���W~4qh�Ǚ锘���f$�Qc{(�Gyp�$�oβ�_��^@F�_qvZ7��̽Ai퉸���ne�q��*�&H�ẑ�@���6�9}+����9�	V\�~Dk;�\]h�t�M(�Ә�(���Y1�Y,}�u/�yoGs����׼׌�6����V�+��ٍ)�d����n�4�F]Q�ͼ��͑�5�/DY�:��z��U�eBt�.��a6V�7������
��k����[m!Wlɶ��4��Q�KE��$4s8�d\lR;/�z}��}�r=�l����B� �߀����׾�r�k�ەq��Br��x�$k�`��{j�DB����@��ӹ�q��T0; Nj����W�.�*L�ޢuoFORl��=)�1�! ��$?t�%Z�0f�^H-��l�7:ҜnO��cA�*�,���No���%����S��k������L]^R93���o\�EfbbkS�S��MO�K�C毗���BY�Lh!�]�Z�3�J���Y�M�+"J�x����<y��>��%���>b&
,�0��a�z�� �ԃE},�pL��9�g%���n�T~���ed"�c,�ma������E-���w�����pM�Es���ҳ��I�HOF՚�\�:�����PkA�6 m厴
sk���评
Ó��=E+�g�tu��O���16Yj_N"�g3��� @�u!����L��+C����m�Z1�u M�P�	��N
t����ŕ���⾴ksb&��*��"��L��*ver�@'k!�ܥC�t�rv�-�DO-�D.�T�O����jA�6Jmq�����ʲeb�s3����3cj:*0P����k�̓��T2�/"'��9ق���|n��&Hä�k�Ż��;a|��a7�����3���d[�z)R�Α�|,s�o;�k����(�da��TG�4Q����uh
aB�G�_N_��!u��oM��x��A/�hw�^^�<@y!dy��`+Nx��q���h#��zM>`��o{K���%ju�.7���4�'�n��C1k~h!=C�㘭����I!duL�#:y����`a~/��H}yW׬Z%g�x�K���-5�~~r��/dz{i�ݔ�eޒj�CR��M���.m���j��Rq(%8ҹ ����T��w3	}��«�ϭv�������!c"��̡An�]a����?�E�ѷ��7�^N�Bm��x7����t�dk0z�����.C��̮Q��$�X�EF�鼥�-X��B��$��?�<#��@�3U�zq"��C樦/ja���áp0���ԶQ�֊�(�ǋ���x_T��T�6��4U�1P=�F��j@��4<L:�?�0���g�����d,Bǖ��9�6j����h�!W�,П���U(���0GWX�l���(��P<5~��$�|h�t�-���ឍk��|����ۀz@��V_�%�Y�>��\�̍P?&�ށJ�m�$;ӕ���Z�Uօ��o�߾�k��Kʴ�r$8o�F�ax�_��GY�m)��W��< Ÿu��n8�/	N���p�s�y�#��>� �H�L��	DH�z=G'��W�:���LW��Bܙ��+G����8O�zij��n	��P-�LՓ�k��q�8.I�)Qp�����g${i�ݦd�⪮9Or-���/Ȑ	fx;Pt�NγԁE7�7��-d/�ӑ��$���{b߃��")�U��ql�1��q���(���F�M��2M��R�+"W�4ڣ�!&(�~��q8�I��]��#�֤i2s2
�K�(��ʀ�w9afV�j�Y!Ni[��@�u}�A�Seyl6��֏�>�������)��LR�h6ɪ�{B!��\�?���[O�ކ��p����p�#��f���u��3tgUTh<<��M�Pc+!Q�I�:w�V�:w�(m�MF�p���.�m����G���p��+s��`TR���3^I��3l &����$a��@_0p��L"�!ƐU��H��Z�g%xfި��6�.M%*�����&�k��;���6��a+���'M�MQhi�Y�j����0����XЀ��I�z�,'ˡޖ5���)��JÑ�h��s1D�2򅘆܄cu[�Yu���5O�_�"�$�0m���.��.Y5y�@9"ҟ����|_-1X �G����҃�Y���T�W���q�3�ŗ��+�0������6Y��-[Qz�n�!�2�;�X����v`�[ϊM�Z�n��XlxVHYEB      e7      a0Q� ��x�d���m�8�"����Hx!T�冭�0}����4�)��S~69	/LD�����ʞ4��[lk4>�?4{a��֓~E�\��U�C�c����=3�&E(gM��n�YIJ���.����82���*s8���`�	�e��el8f@