XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��*5'�%ҵ� ��n�\���$,YYO��0PgK`�����xaܺ�U�l>qZ�ʵ��I�={��5�%ʬ'OB&�Bl�	��E���É.����7�7nB�1m�%��KK��I��V�,5�G����3�=���mn�r}n2ﻇ]�/��1�^\�{Ϩz�2�4�w�c�G+�Y�t�Tbn�F귩 �*} X��@�ixD:�����ŵ4�I\�� <8���&�#J"��{1{��W������Ϟ͝��ת���$qM��=�X�8��>��_G��M���]�0��m��S��eX�1���0?�C ~�Mm2�+넱��Y��t�O�O��Ɠ��%�\��Y�g!��	q�8���P�PL�2iogHg`���́�Uѥ���]ֶ�����|�2<%�3��޶u��0��G�ڈ����oGYǃܾ=P�Z�0!��;�4��_�d'����뮘�4��50��<�����(�k�_����@�3ͻ�#=���C=��\c���ϔ�n��R� ��1|v%�+{��랫�S6|�v0�!�!j��յj��M�,u�>5A�߳`��������x���\�+�)X]�L��ߏƔ��|N|K�-�t�U�?/$���>�p�^�2/��itR�h鲁���m�_���A�Q�k�C�Sσ>%{3O6?#�Z������C��
 ���l^�����
�[�r�+�3����{K�ۄ��"G�oM*���U:�Qb�Abc0`XlxVHYEB    fa00    2560ж��P�Vx�Źп{�v��맼��� 7���Q&s?�L�����W�N�+��?��cݸy��*pw��;ZL��z�JX\�7�YC"���q鸩��vm������P�*<]I���z���_�B��?�"��M��;d��o/�D�њx�H��y��$;��2w?.� �YܪE�YG��7 �gm�0� >o��"��\��;�\o�98!��օ��YX�%`���+f��C����*���2�N�	�׹ˏ��\�;��_sTY����q)#�y��LF��l
�`��2l�t����Ykm7�.17�_%$����R��*���Q��^�xu��#�OSe��3�1%xw,�Ɍ)�	GN2}ҤV �!v.N�e���\����')�9\�{c4�/�ݢ�j>u��=�|mp�9��34�-%ce^�R���Z5��ή�@�I���=�[�n�-"�v�����S)ob��y���o�R&�'�F-B��m��(q�[�U�I��-�,B����-�}�9jr� �z$�z���������e��Z�	K��� �@��z :��Щ\�ߨa���7uFv�j�Ѩ��@]�f��7	�DwzT�s��Y(�0���R��p��-�Y>�ύ-�L�$ �w��E�I�e�B����#XI��O%�� '�]��o���j���|N}1i��!���,�V�J{ai+��Gh8�x�⣞<F4;K�K��Ndpl�� �|��e������_��j��#'B�к1�S�_\6�����<��>����
5�BT(4h�r�q�d�è�|�>�����R�j��`Au�_RR�ٵ:��򨹠���d�8tx@J�2Bfd-��u�~<�l�	7���������Pu���N�x�*�ր-;r���֥N���1����-zO�K��UQ�ɡs���X�
)�����)�R>,�tnm��꫽翜þv�r#�5K<��AR�~�����
�3n#�:��b(��F��v�[�T%Br�ȉ��^�O��a-cg��[s�EU��'���'������&�$
%����b"G>�,?\�r�Ǐl&[�g�H漁��
�c�G�E9���Dn����ǧ,�p��X��T�~�_�"���\{�@~?��j��X��p�v��*��\�o���a���oU�t��6�a���S1�g���	!7�i�R�P��=�~/ܘ|�4:]2\vPm��:��\M�M�u�9��G�"X�e&>?b�j�͟^�%ð[˵�۲6���'tNh��li�b ���B��]�em�	?��"kw�D�'y:>	~����{�����,��tU�g0DpD`X���Y�{�����1%���!��B��|���c�>5����ȨLt81f4�������N�f���\��>�ŷ�`sga�QW��lj:�#�z2^�Y,6"�Ʉ�$�'�#���������8Z_���i�� ���w��ڿ#���q�/g���X�K]�%*��ei���F��~xk�Q�
'�x�����Q��r�𸜰�o'-ޜY�V'F�ag[ڪ��uɭ�}(r�OA�	�2��>���wz'�ݾ8n�Jj�ÞF;�y�3��2
_�����W�p��m<<N	�-u��cH�ֻ� L��Zͻ�_Ǌf�=��.H��?��=�o� ����z��8�V�q8���L�4 ~�k���A5[f
jA�n��؂��������F���M�9��R�+7�!���K���A����ɠ��,Fx!��G���XAܛ��>77�>4Qݥ��:�k˝�5~�k�֠�v�r��6���&����M]�>�i�_�B���LS�ß��|_Z���l.��yr�&'J���/3b��j�=}~$6�}A��Y��q��h(�jx�x$���+���)?��P��'��n����Y��V��%�\z@t�S^�K]}NԌac����W��'�ds�3���~s�8E��ak���r��N.�|�Di=3K"�K��C�?e�f�(#D�jt�$���w$rnC韃��Ѐm��Y˞��^���n�����lu��LpW�Ծ"��р@E�R��y��4e0�Q������G��X���0t���T�!��\��ܝ=����f�ج�|�s$���%'��!��H�hv�OK B�L�o��Czk0c��ϨC:J��JF���Sq��Sy�kK�]�S� Z��KUϣ�+(��N�;O/PI��luu���dt���l���st1 iKK��MԻZ �`�	]~��Q$<�|��v/�gv�W��آ4����I����z�i
�p������C���]IS���%��a{��̿�L/��Tp�qs���m��h���f��� ��brO��#-&e�@s��,��l�M=�xdږ�NhQ�i�z�`��y�Է���蚋�2�̞�Ol��ܭIC�6ر��ӵ[n���2����.騵����.1�_;]b�(�=7�F��YV��"��M��!�u�~�x������L=�!zqr&�aS����G��(H�q��".�{sߟ���6x��`Ķ�Զ�b=&;����A��`�֕
��M%�2�;/8g�@x= �1�;x��#Kg ǎk<�T�V��UaC\��yG�= gR��b �Ix&LAnx_J��>L7Iɨ�r�vpU�� �tTN{��w�/xVs�'3Ic2ws� .y����R :�Q2O��>v?��wW����!X���x�܋՛u߲��ɪ. �	�<���>���i�ZI��t���{t��\����8פ=��y����9��W�d�Jm�[&�~��$ǝr@���&�ɇ�*],C��:o�_�c��8Q�,��ʚ������5:����,��s�H�"���m��1U�s�pឃ*���
�!=~�A ��獯VV�鬺P�Ʀ�k���s9U�x���Ж�B�z�g�~쀋�+P�+�Iz�^	�׺�I��I�Gh�XB���� ��F�S(2�2$����pX���Wp���9�&0�z��:��f�1��#�1J6�k�O�iS�M^�Lx?k��8e\B7�aws3�p���-��j�Wq����}Q=:eH`���*7�	���r:uG���eM҃�Ƣa���j�"�,�0���<��Ǹ�Ό"#�����>�Eq�A|�ˋ�l�kj���mr���nS����sF�=J?�f��5/W��7����t���&�޺�'q�}=<d���$q�{B��gn���o'J_���:"�2%K�h���by�d�����	����&cG4��y���>������Ʊ`�9���օ�Rp�u�� �ݮɧ[���Y?�Ch6�^WX�Ȓ[�4�bF���Y�����~7��O X�?��.��@v_�G\�g~s����*�i��`����.i��� x?Vz�+��v�s�.K���ɟ���-�Hs��@��ٚ��HC7�����إ)#��+�X%�l��D�
G��.�oM5����^�v|�R�X�����O5��{��8�"����Zb�@#�3��
],	@KD�M|Tm ���Y#Kj~)�?9�Ak��6?�X�/|[w^�t��'z������*�<��;t���]+���Β./Q֏rV��j"46�<��B�����������>@Dg��6;!���̢!��t;I���|����)��tÅJ�č���>�~�dH��U��C#��ON�;����e����EY^��g )���$
���CM�9���)�R�vY�R4��֎9�[)z��Mh`9D���w���Ȧ���@ӵ"%`m2�����ǊG�TIs���c�~g�)C�5	 �:�4����1ߤ�t��L��;�����{�·@�p9�|,�Ҵ3d�d�v�|���x�#1����p ?4�,t5D�d��~mJ�5~A���W���������%�J�̂��\�gY��٭�{n�1X� �z�/�#���w�_�������+�Rk<�+�t�z�&n��&���x�=�	�?��/�i��n��mY���%5��X�k�L��8���k����=#F~��{Ǟ�8��~A��w�V��4+D��)�����q�Y�J2t�@��ͩ�va�\<1���㐥=�l���9��qG�m�f_鎚���]�1��!묄�XkT�iX�����@F���*�o�,����<�]�y�H�GL���%W>��pl����z�U��L������c���^��R�0�v�]�xMCn�CL:d�<�[L��ζ��Lv
�j��_u�7?���h��4�m�izQ �}�Khd
�aT��TH��_,C����O�y�R����ἲ�5��H�-^=R�TD����l>��!ō`I ���zLd�r��d٤G����ܗ����-);zfK�2L�b�x�}S���Oekʈ��&���|o5�L�5�%Ǵ� _KLb<'�E#;�G_-p}�����\�mu/�#�^(�RIӉ&��P�rE<ڐ���%�+��9�� 3��/�V8�n��.m&5Z$Vj[<��=b�����<)*�(k�ƽ��:+��T����v����/ļu����P	��$���?4W6Ƶ�~S��@�"�1[��Y�����!�c ��-àmk����=�.���Y�g�"C���9s���Y�o�ڃ<sT�3�@�q D�;;�j�"p"*푝cG���g~h��p.�����L����?�@��_5<�� 8r���9�WcǨ����*d��"���Ƨ�g�z��^f��#Z��}Lϗ�K ��8ʥ̗nO}+W���4w�`�*��i(�.n�gsj�
~le
h�VO�T�Q!V�[�/:B~�>N�[qo�C�4ãI�A����)�n�P3�NFR~��-;�g�,�V���g@���A�wP�5�Ho:���Q���\��G�~�e{&���M(���������%[)����g��oa�f���q���c��RW{)0��j�/:>�K��]����|���t�Mf}V)�xY�#B��?M�����V���7�[fO���vnǼ���H��]�{5��ܱ ']��e��J,qWkֽO�)�[�}#��Z'���f�6��g�y�f���2������5�(M۸��>��抙�B�o�^3`��z�@*Ε8�X�>F2�g
~�v�w���'����4�]X�6�Vb�ŸAا��y�-I�DV��jN�(�Æ2��b��j+�~�2'Iָ�s��j���!�v|Cgk�~	~�^�E�l�d��R�U�X�԰��Y'��=�ڍ�5h�8�f��C�7��*5w�F�yX��<"�LB�t������X�JL[c��O����)a�걺�H-zd��	#aS��:��e/��y\3]�r>g�z=���Պ��T�T�Ix�a%������N����Ћg,�D[��|��I�RrL�gn�AoQj�wܱ��;&�^�($�M¸��+���l�_�YS��ĳa�s�y���hٗ�PV�'����ƞ��v�<g	Y1�
;c�Z�7�}o���ފMF��pA=�d��/*�oj6B�(x`�Ҳ�4���3Gի��%c(�Ci�̤�+�0�1m��T�W{��~�i�M�K�ק���͏�)E>�xo �_E(g_��,Q�=@�*e���^��1q��&m�_dk��֌O;:���t�^jb�_"�))!��f����>�E{�o�
L���3���
�K'Y��޳230ح۠GE0�OE>��?��	DQ��K�H똩���M<�O6P���U+�{Q�ٳ�3YCLY7E��{?/�Ou�r,��t��,��?1�l��R����E?�#�����H���q�T[x�ʕ��*!�K��m��Oΰ��W�61s+k�U:����tG�K�3#su�H�!�����dW�vZ����9cplv�^/%�Qh���竦�z�z�X�c�����nE���=�U�̖sJ�*okB�DD��/��@�`es�]n����
�0����A(������r��R9��l�*Z+aJ!/@�˝3�ٙP�f��R�H�R6`���MS�k_t�?'w>mě��{�?�!4�T�H�Cӓ�w��C�sL��k:q�Vu1!e�.=� �H�>��4�Q/<jk�'b�]9�C���k���'˒T�8.��p֢l�惥]�Gl��@��R�p��{py[�$�C�~ |g�n�����=I����=,^��w>�k�&?#�>��?��s�P2f��O|�������B�N����oZE������m��!�b��vXL}�"�(H�c�|�Q�?[d���k�䉝�a~j=�t��mL�0?.?�^���p�����w�Ht�^칩8�Z�\�:���i(l���e~��V�<�U� �_-�dJ'��N��	����ƛ�V���đ�6U�G�y#�E�p�&K�<I7�i���飺���k-E=��`�9�P$Ǧ')�3(��c82����aգ5���㌧w;�.t��N�x�����;��7��A������AȞ=ZEw�׷/*X(r-c
JI�V�.<T6+�*{���x�LL A�|o%R��Tk�P�]�DiP�L������|\�w���Y�a>,?zR�DAeZ��B ��Co��=�|y������������6���ݙ�����-:�/4�و�jR�k��/	��Ak��w��^ɻAb��L��:�ݠ�#W��\�*25�,p���=�d9��y_۾|��'Q@L�Jd�i�޷p��)W��HLfʆ����hG<�M�9��mg�^F��� /���=���V�%���� !����PD�H���	S��%��Y��O5���Z�A{Ts�>�Ϸ9�f�ܗ}Dˍe�`
z�0����9Լ�$H�D�Z�q��R�~��p���D*#
q���<�:�G�>��ȸ�;{�����o\hs�d�\w�0ۺ�1{���hU�������b��2���t;u�=�GC���^��o��<\�4n`^F)6F2_�_���z�4�K���;����X�U$�<�y.��B�"����-:���s�����\�/�pf���d��08�N�;2ѫ[m�e��(&u�u ۵Q�\Zy���P��/W�b�r⇗��^!�:»��	�麃q��dC-�ϩ��~�����>�"[W.��XXOCJߟJ$%c�k���@��ڀ������J󤐦^��E�r���t��d ���>UG�`�O{�ZB!�)	�V�s���D$����@�����ݝ�ߋ�eE �eQ��F�mr'��7x1���fk���<�(�E�;�a���,ウ�y�*�IG��z�� ���5U�Ǎ\��wS��X��]��(�G~�>#�16���϶, ��z�wlfxi�L��<\i,�*1��1i�a��S@J��x�1�$n��q�rh�
��j���"�A��5��ܼ�Y�쐼s�.�i���>��d�KH�Z4��o�C�b6�3;A�빇�$��渧�W��NQg�#��_1H�Ɔ�ʝ�k|�֟�6��e�Z��.���G���޵.+�Ǔ�.�k�5C��0�oݗ��o��%��6/�BF�φ�iٿ�Tq�[Q6/��Ӎ���4ڭ������$B�8V{���#��}��
Cts[���T�Q8�i��Fx?Nctv]��ˈ�P�@[�<LL
��m�*�������(��5��L������{�F���E�l\����4׺��RK���Rk�!����k�$P{��F�]G�YA�����~T̗eq�.�h��*�|U���^^����6)T�s�DoV
c��ݐLF�~���TT�xށ�S�Bڂ��Q.e�ꬁ
�v�"_�	gה׊�Q��^*�;l���n�tV%�¹G<�ya)��*4:�nJ�qO�t�2p�QM�Ҋ��Yꬢ��󨣒`ƣ�.mƎ-A��V*)���B��E����F�ǟ��5o�5~i�1���ؘ���!$�	X�o��ۄ��������/�z+�&lYT��*�� ��sЃД��g��O��(cBl����o�=煰Y�Z���la~J�G�>M��F��6g��������J� ������TR�;xl���#�^�ÃGTn���2Q���ѡxX)���	Mb�1b�X:���%��XAQ9���[@mT*�[er1`��A��=�r�!�!%���@*���&x�_Iue2��8`y�G*:��MRbo����z6�����%_цYЩ����h]`��<���#�rCH�lV�-q�Y�~�2W�DMd_��<��F��Ơ�n�uU�MV�~|���WY]�T�@b����z�e!!�nm���S��\����|;j��U�[~ꠥ�g$����M!�*���*�� ��^���\��"T�Gϟ�k��ϟz�[l�����oD��9Hx�q�V�6�=��LǓ��װ�� ���1;R�[4�1���qɴ�̔f�K>�������&��[�)���R���+)$�.���'����ѐB�^`p��Ş�B�J���	Y��#�boӄ!��pq?����������Q���$m�,�Z����	ȥ��l0�&���
�gG���Р@���ht����˫F�����)�!P����+|�X�G&�()w�e�H1��,�<N!�M�E���n�l�r"$s ~�G,�� �:�7�z��Q�O�����
hq:�<$�&�
��Z#ig4ݒ��Ԧ�Cb4��i��dU��҄�^P���� �I�ɿQ��*sۑ��-M���*�vg��=�<�P7+��!>��X��
�g�~1�ֲ�C?[*�A�]�z����;#�:��-fX����b!`a)�u:�c4y���+z��}o�]�Z�ٵ�OA�NIe��2�p$-�.�n��'3�M~r��%��/��cu���H���qu���:R{.��)9��[�S�R��Hά y{/�Ȩ�<S@��t�˗�U�z��Zza��0�6��z�1E>�$��oe�"�l�<6F�m�p������l�a���'g�A.�����q`��}����I�e��.0uIQF-�S|C�K\�V��z���+V��Far��>!�}�ӻڮ9b�DH�k���x�Z��}Ey�=�pk1�5�@��;H#Q�D�xi�Sl��("ȓ�$%@�}t��������j� >�o�P�-T�� X�|�<2YL����0�a>�3�H��.G��0�B�8�%�@�U1�MfIX�p�%V%?�?P.$���}F��A���׏-x������P�
��:�S9�@��e�t�:Y���ix]�G�zp.s�c�V�_���ʯ�cA���=-(`����s��^�m����C9iY��}d7�ٙ�S ��o�4��a
b�V坦ͬ��Ep�E�e*����rc.h����Λ`֡v_�J
rn��]��[XlxVHYEB    fa00    14b0-:.x}���-�z7����oPq �HY�~��rV��w[͙�<� ���REB%n���i��w���ݦ��̗��P�)�<��؉�*��Ο�9=M�>���|S�P�Jn� �5�#[N9ˑ@�o?���sѣ���gm� n��9�ڟ�l݌��8)՘5��/��?�+�=��^�W�Q�ۖx����W�dƾ��'�	z2x�0�`?q������!0��a�~�4��Ti�0O�K��=(���o�<�_v
�3ߐ��e��9/�˾`E3�sJu'D�����F.�_��FK�d�Q�]?W�qOᥳ�af�Mxl�c
���n��'��&m���?L�����i��ܰ���r� �'�~��ڨ K����o�嘰�����!ؘH)�4L[��щd.�`v��|XY��Ŗ����d�c������!��o�{m���q�G��/�]/��
�T�'�_5�Z��9�v]��8ґ���AA���i
�=�eYR�B����rGsfO�c CD���]��K��T��5C?�Q��s-(�
��.4g�t5��U��O.��b����rn�A$%ae���[�N4�ge���N��,�q��k�������{k+^���Ey�KH|g�2�H�8�mb�IG��z�֒�']l����C;Tˉ!,�V��Ɇ������'jPPv�݁ ���&l1�l�� �V�_)SD�I�F�E��\�����P�E�tI�ZJ�����XaRDh*h骭��[0)�'b��/�B34�Qcu_(Y��S#������*�g�3lޙ	?5чwK���M��q�����;c���]Vae٭�QwE�}S��,��CyUi�o<�1�~z�ר��,1��]�K�C3G��tw7�C������5J�yr&��G@�)H����1>�c�8.h�I�~͜��Mn[��M{����G^�fus�*��N7�ԝ�Mr�3����XF�(�m8g�2sJ"#2B��TL �-GK)F�'�v�KXyV��i��E{�*�p�����af�=�3�i�AXj6��}+�8:\��l��U1"&�_PJ�#�}Sj�x�62)3E@V����cqn��_��#�TތSzT@*����T���Za$�,-,����,ځ�]p�v@<�q߱�ƨ���n3&�k�aQ�v�-��q3�j6A���JUȀ� ��ImY���)�0H����oqC��A�@�ikkɅ�2J�:R��U3�U��x��#�9;���N��A�>��nع|s�Q�A���L�ʵ�k�ن��[�����ic*�iR����+?�ea�f+*2�:}W�|-�;�Ԭ.3��(�L�gVѣc�B�)�!a�)���,���SI�<c��|*�:f�>p������[�F)�@n|�da���#�f�{ǔk���1o�̢��*��3��{#�X��iW�.�d�L��:L"ŕ%��1PF��6Y�jy�p�����e�%��颹�ulw�I�0�e1{���'�ٜeoc�}�z�g��r�ʜ�3�]:w�������\�^t����34޲���*%��C}D͠)��p\���L"F[��(�7{C	��L�U���� sL�j^�혏>!��5��2~�@�Q<��|@���'�0�<	d��TY+��`5`%Y�]r���'�<��� ']�	5L�S׍}Y�"M�#g ���D(�^;��0�%$�:�|��|5����HY����$�N�A
V7q�A�/��*C���~��7i#\JPJ��Ka�VD:� ��ZA6�^�L�_C�Ňb�.1��a"jB]�N�0��y��κ�@��lb��P�3 -ݠ�tj��o����b:�3t�L���^��)rNۚ���
|� �	�
ݭx:5
����'+7�(<��>5˩����p�I��X"�����
�h�՗0�ߠ�L?�Ag�^MЩ���6 DFc�e�V=#��=���C�L��_ȃV(`U��[qG�{�|�_:
"��\�F�p�i��j��j�P;N/'U#���Z����LW1��Z$��m���0|�Q�ڿ�B@�R�p&�8�������CPe�f=�gP�w�h��{㔎T�j{��x�6���n&�ҽ�Pc�,���ٵ	��V��p ➶
}K���oq#��e�T]�h8��[����z��H�x�YKs�* CU�ړ1�Y�"{5������0���=1WS�Aw�O
@W��;�����-���X܋!: ˜��M��E�<nv`�|Ddt&,|��/p�b��`�lƣ���`�5y���QVTr����^m��q�y���/��`� ���.}�2Gu3�ҵL��8��J�^?�ȅ�j�0��AW֏�Ċ'������A��Wj��٘_Ce[�T
۵\�E����n��?�)0u���lѸ�>�"�{�0Z9�akb��nw�Aw�US�v�<J��_��ƥظ�\�\��S�����(�a?��U1v�����w�*Z|��~wXP���p��.}L��C�q�-m�$~J�>vi�k��T�8Jm�`����x8(�St�~8R�7�,c�Q���,!u��m��e�G�����o�HfK(�W7���/u�����Ai�J�c��謿�������uj#a�</j9�>b�}���;x3у#��<����I��$��.,R�	�U�?��<��Z��l1���_�Gr\6νx7)����/��&Vu����h�1�Yyv��q�v]=]�b��'���q�5����E&��xH�>3��{�Qf�/�05�Vݯ+��x�9F!��I�?��-��{�`�RR/�+T��l�y��ԑ����#��r�|�Nr�\�z�I�" Ư+�e;�@��;J0����y}����0�UA CN��7�
��j{9-qnk�c7���C�:����֖|_�J�y��4�"�.��U�G>� �	K��Z�a����i����ڰkk�dGf�9"V}����?�s�Y��P'.tu!�H������f�92" [7�WF8�ij��y��l��D]J�
�� ��F9���S�:t��Z�A8!���l�V�#�1��� [���;���"�ei����6	�����@�-�v<�r$��V�`���z!;u�5�\q~�7	�!Me/���j_��LF$_�i)��p��0����ߊ���d��MC9�]?gw���<���:��g�_v���h����Z�;���\.���l��&_.<���ܫ�h)��;g��ۈyp�$�x�!l���?�Ҋ\��w�$�>+�0܁����,a �A�0O�H\5�@���`Kq��bf����~{��{��C�̚��hH#òY���M����pMᏰ�pX�1�����_�#�q�H��c7r��BX( �|�z;G��6<,��$$�k� �t�u^m��&7��!9�쩟<�K��7�`��Imlµ��;���b呼����o����,�^pzk���ڮf���P���s�B�!w���}4�*AB@������/�f��l�`�2F�,dj=�r�%D璵�,s+�D��p��3�󠔄��M4iBH�Ů�,KD��������p`���g�C��%n��4e����#>�J�|��_9~�:Ao��l�|B��rx�J):\���5�# S�V�fC��5�y�k����&nĪ0�h;	y���U#���'r��lCB�phIDA~�V�>V�^D��/{��
	��n�;yM��FGF��խ�J������V��[_y� |�4�e�ɱ�ӕ)�U�sZ�7�L]�9�ڈ�n�wT�(�7f�r��T]��zs� �D?�q���LHs�N��|5�C��a:�f�ŹU����.Q�\�t�O7ؕ�� a���~�9��w]���؞U3xf^��x�����z��ݝ�Ҿ�/ōag��}�����N�T��U�$�Փ�0��BJhd���Ѥ��h�^���eV�$<Su�J!�3�,y£��4�U@�[��>&�Q(=I��="0�h��Z�ts�ɛ����;�+#p�D3���g�t�T�}��m;5��f�����'��NݠYv4?IE(%]9�Q�� ��XR�<���XIb�yJ��G�z'{�<(��}\�{��دQ2Z�2޽К�,~��΢��p[ =��aGE���R��D8C��`2;��򦣪�2�ȯi�Y.����J$}�&��y�՟�E��M�~�Ѱ*fl�S���C�s�o��;{U��h�L�@�eb�K��[	�kxM\R)��FJK���$�����k�,oI���'�~��ѠH,����ග�������d�1RϜ$��sW��N��jq���d(qe�:7�M[봺����'���7��:�8e���]�L�@̀� ��:��0�@�큕z�Vi}E�t:��~�������;�ۨ،�M+C��ά���g�/_Cߦ>&���[`��,qvп��o��zgS݈�@���z����dbY�]����J����#j�D�1`�q�l�5����	����1�A�N��ݻS����ˌcf��D(V�wv�;}��2ժ�W�1췆�(E1�ee�wGo�{������� 1�M�:�+!�jT	��r���
�E;S����㽂U�,�G�)^
a��L���k�Gk$釆c�}Q.~��T6p����#�/ʤ5��1C�#�m���ĪC�ֽ�h(���/���=�"gB��=����'Z^kux����c�o�>�T���^����'O'݄tFp���?�	|�,g�%J�ƫ�m�:���o-bm� ��xN}/�`{WCO��ρ��U��wIǺ����1�-8ݯ*f57n�G1�ޘ�::GO	`�u[��YV�� 1>��0�R�[0h.�5g҇VrWn�!��i�Uf$�rHd�0rm&ۊ$2�k7���`���-����21"����Q���m����{�H�� �	��+�zFG��z@>��L�¥}FY"��⺃[�d�A�+�ɽ�'?��j#���/g�v^,�\��*����\��'C�6P�/\�l0/��3;����1�uէ�PN+N.& ���9O���X/(�2��] 2F�5[M�tr�pa ҝy(�F�I��>չ�x�tؑ��i-�ꉑr���+�Aq�p�	�������s<�c����Ў+�^�/Z�A�W���r���T���3�1B�5��]�֯0��II-�(MS�P�Q��<�C�)	g/�wx�Q���D���r�XlxVHYEB    fa00    1880�'QG�י�5��^�Ë�����b�O��s�}I*�X�t�h/���=v6[/��8��%ܭn����;�W�)���i����j�yp�(C�6 ��`p��l�~>6�D\��4�W��k�Ōez���Z��t�P	��{��F��h�v�	0R rx�+�ֆ>WU`�3"mIO�լ:�.���J(_L׊>+�����c�/!�j��ӄL�n�NZ�>;�T@7iHdw6���DS�٭O5�[���1�-+�p6�I�vpҙ�ax�����n�����l��L���f�WZ�z�
/�Hj�T"tx(�F��1���VN���IAO|��
G��^	�������!�Fc��U��Ҙ����\'G��s8���r�V0�*��\Ɖ�����ꌚ���ƙ3���.���)=Wq�svlx�M۫���֍�(�w��K-�iM>"���ܶ1s�n�z�(;d�y����:�!��t�}��y�NmXM������~�f�70����X�EO��o$��\u\Y�Q+ i」�. ��Nse
�5���}0�_d�(F�w�.N�VJ��b�c6�:���g�4NB3�n}�~^��).%jE�p�ʊ!D�� �^�zu&X/�>a>TUT��l�E
�L�C�
���Xa��'f�ꔉ�T�\�z�R*z�!B[us��蕍ș�� ���o�v�/�F���m3�GU&��*���c5}BwR`��&�DF��zT-M�"(�e,�}
�e���C�u�j�G���
�騥[�{��	xC��������ZA �1�MΣhJ>�UzC�P��eL%)��}FZk�lk-�k�.Q��"��~'տjj6}?���({4���:����.$]���z��Y���b_��=K]=Kc-�~�vڞ���g�K�F�=��*d�o_�nv��G-K`���9��|\|Z�ؠ¿c8+��g�A�{�upqؙ1���:/0��F��������	H����1if~��C��[Y�NG̭&l�����]��q�Dq����G��S�m���*��(Q���q 	�7z�3�@�����+#���U��Z������J�l�k��X��P��&��V6f�|��k-��/͙25~мp�ѥFA������G��Q?c ��Y�%���f�B�v}t�P,�]����jè�B��@?��f�CP���4uC�W�p��˭�	q�Ss��Q����Rn�D|5��6��%N(�4.��̎I�73{h�
u�ʁ����/�Ȁ�n�N��G�G���(�6~-��8��Q-��	��FT�[�Nva��81��٣m�<�v1������77y|�H�^����Ґ�k��ɴB]��@@!��+M��<6<�Y�=��S�6ɣ|���_�b$��p�:���^2�3K��Η�b��TV_����Ҩ��\s͞��(5zf���b8ߜova.�V�C>t�Q_�5'Ԩ�v ��dc�K�&��#��_n�:�C�_`�ɧ�����,du�b�a�wd����j�ʉns$��rl2}���wCp8����g�#'Z��b�b�`�ӟ��J�����&w�(N��UQ*�D�*dH�hn�l�荘2��n�ӦDb���tP4��������cmh�&�R׃��E��;ۮ���A����z55?M���Dk��A������}�&��S�Iy�+Te�u��O� �oO�qK���0$5 �����x,L҇Y�q�P�k6��<�u��.����9�	�K�S��xۢ��(�Ã�9����v����){�:k?�E�񃒠�4琡vU� ��wX��}���RD��#^���S*����Qa�1�r&��Ǚ��Dleh�"LS�Ѵ��ǢĄ��ρ-L��a��ÿx/��R����# P�&����Te�Dr����g�鹦"<�Z���^ $�6�r��zE̱ruOK��s7�?qN>�j��s�n}]�J:O�϶??~).���r��K@�u�(J����#y������.���Ld��,�HY��r
b��oi��4���f����јX_UR�t��/�p&�g�t>��%iC$��Ϣ�fl6Mv�nH���OV��в'$~@�a���eـFDlq���"���h4f����U^GH�aȓ����S7�u��~{q��a���������Ѳ��_��"�����%�Ћvgg��6�e.�-oA��c��5�	�ƻ	r�|dTj�+��J6��ُ���Y�iO`m&ƒu����y:�a�:���L><�h��s�3!��/2y���񯵫��=��\'�+����\��*�R�KG��T O0��K|~_;tf�k���y/r]��&s;�E"3��>��5�T��Zxě����E*G�G�$78� Kw1�<'ʩS2W5b��ЂKX�G�Ve�&�|o��K�]�o%���|J��T]��A��{	M��~�Hv��I���l����w��]�h��%���(�!Z�
93�<����3l�ۙ������W`p�G�Cg���O�L�-����K�R����1�(T�j��Say��nS���h	�� �
o�T�]'��8I��^(K��lX�P�?`P��Y4S�>a��uD~1e���iY	t��%�|�=gx�%̯>�#`�'�6�w&P�k��+N�!H��,'d�{�} ��"�:]Q;nSB(��)3w�����)���u��txǻ��Ǜ��3�zp'����F� �J#��5�\
�d"�\������7>a����
��z9�$��JB��^��Ѫ�HA(H �� HSCq'���<�C�������MEH�%�N�,���y����EѸ 4����%���<�D8��~.���sͣꍾW��z��,'�U�#�uQ?�iw�:װIy"���M��)Y��셿2n��� D�m��J��㦕hϞ��M*�gф�r���@�B��F��,���lŜ#���[5+'R�~G}A����W	Ψh���I����ώ��fu;3�_��+�6�L����dE�%�#7�K�Go^���ޢ�����������zŚ�3� c$����<�(�T��y<�+�Sj'����ҧ1��d���Pi-��=���̨�}�)[(>�n'������
��@ږ$3�d5�l�*�W��6,�2��i^��Ym�e$<��R��=�������F�V�P-n�~)��H���U&˂2�W7��'o��y���}#f\gl���C!̋J9d�8l�t�6�hH�!���C�U� 0����R�$ �r�H<�AV�yg�F��m��X-����K	�P���3))���7�TGg�J��zm�J6�u;w�)PF,ˮ��g�R��A[5M �@w�9˓�8��N���>�ΠN�� ��3��<�g]긆/sd��c�Ż�y\Y�R���C��)�K�;�{8�8�z�S�5f�#�e+!��3���Ňy���|;x{g�y�y>�t��s&� ?	�~�[�/{v<�����C44������Ͼx@���J�M��2N�66��ٛ����R�*r���J
�7�B��a��W�@-iy�k���u�g�u��^��G�k��W���� ���D*C�Qz=�>���5���f��FN���Z��s��4��I�ӥ�C�oz��Cs��^�������<��5�t��2S�����8�%���sޛ���EL�x�U��Y�3%NG�oLӫ��85*�Nr}�*�'��/x(;��#�<�-h��ù�$�PF�&�XTT�s�p'.��d�/}��h��!c�j*�����Z�a�Oj8=/�X
����0�ݸm@?Rs9!x�8�	JH����$y��)���O~j��Y���8�\�#h������;����列���ѱ�Y&YK�`yeuu�ӳ�{/s��?1��g���w�H��@J�T< D=� ���fǤ��ڱ��i�4r�p�4,S,~���S��������K�ZQ�Խ��r%YZA��ʏg ��c���E��ξ�v�Ջ����E���� ,]y�?(��o�����1yC�il��мR*R��M@�����<�+���=j'[w���aIQ[�Ɨ~�ܘf�v��Nޑ\s��?�V��!��Y�y�1��7��M*��ח��ۥ���NG�P+t���NH�sX7���s�ɞgX��cِ~Va��K3%q��RbSV����оi�.��Oҩ�X��Kr[b��	�Ү���X�RĴD{����P�U�ɏoU<2B52���Al�:�,U��p�{:�f������|Z��'�gS_A��t�u���29e�3��y^!!����=�%7�A���Ek�XS��^�Z��D�MY���%�Po���d;\qDʋ�-����{�s��<���#��%F��4���Y�)Q�IK��](L<��KaN������^
N�Rn��H?�y�����iL���8���*���pϢ�j�H�W��c"��T��om����'0��kY8��.��-�B$��q懑��H�řZ��k4�=��Ҏ�{n�-���[`At��:
e���ԙ}ޛ��o�MC\<����(��&K��b;�� Y�vF6�����4�LZ�jc$
���]�1��7�>3T��m2c^#|	��7�H���H�ج�����)�D����\/�
\wͽ@�>,]*�	ȣH�E�0:Z�D�Ď�O�� %�('�b��&���� XIsg��מ9'ak��o'>h04nJ ��|(A�)-�4�n�@²˵���r}��Z"ϴ�@�+h����ԇ�{WT�����c�j����{�Ug�1p剹�4�z�m�/�u����!�u�R2������{����˰����q�fj��B�ww�	�����w��]*��^�	��iZ����H�j���ݰ�̨����gF e}�O�KۘX���e]��\EvR=��rF�Us��f�?hV�_3򒃑>�	�2E��K�N�O5z��7��2�w�[�fU�`�Ğ���<ÑP��V���	��~P@���F�f��M>�k�4a���*1��"�V����L���ß�op�K���6O���zV˕tB��xGɅ2��eG*�Ϳ9d�-N�.�,ɦw�q٤,��&���Wu�u����z/�nԬa�O����O��%�&���w(ګ�"�D@.|By�I���%B��:��`���5���T�1Ri�O�z8_��k?�����G����F��Y�B�C���&`�%d���dF��g2�a���!{���s1E&�)��6t�O��Ȗn �:&���8��b3����y=�G�0lvxPz����U<�>���=b?��+���v���pC9�x+)�Ln�FGu�e0j�!���5�ԏ�o|��'^�z�� ���8Q�J���H�7�%{3�n�5]n<�t��0��-��P�'�h�n^��N�$�����-��	�D%����J���%�W)[�ňW8��`�ti������o��})�=�*��1�H��3���$o+��ߖ�%yJfX�����"$b�/?���/뫩����B��>�������z�?#yIv������{��� IK���H�a?~x¦�-�="Ẉ(��ߋ�������#���!���d������tJ5VΜ{w^7��M���(�'��[��J \�K��Rfx�	FBL���D��A�@���)w��+��V���_[�Re1�A�6I27���:|��U�Z�pX��d����pm^ �y�����X{0*^3=e2^R�.�pH�jF�����a����V�٫�q��a;�2�9��z�ƌ ��)�o�R�ì��e�7׉�h �����V���\�.�>����B[Z�K�I�Z�&:G��/Xϧ}�8�/��AL�qກ<Ϯ�/���8\����9�@}�P���g=���sH��~s����/���(O�Z'B1ˈ�	�1<�+�]u�q�#��b]�R]!t@v1Ȣ9pCHZΓP�f�=�L?k��Go� )'��Lo,$A-$?@�F���u�M'����SZ�=$0�v��|�� ��;|��Vvc5_.:[$_B\��Lߡ��7�7���ޤ�0����W���.�Z$M8w�B����G�/ڑE��G���7�����M8�� ��XlxVHYEB    fa00    1910Ի5�(
f�$?�zƀ���v�┘H��r�nq�[(�ܻYz��d)�aTM�˂ծ[X]���ʰ9��mn�����*�{������B�.�Kd�_3�I�Wc�ǌ�������d��{����Ĵ�<x�2h��<E�-I4?R�=E����~��UO�WS3�P5�MZ�ev9��D�������Q˫���۷�)C�3UΪ
�/�`��V*��nU=H���)=��Ɏ}��4y���O��r..�ѐ3 u�/��$E"8梲��ztu�ُo�u��K�wĠ��-E��;F��kP���&_������ǢsfFLCl��&p�#g�Ӿ�'��ǝ��#sI�7����f���I��^HFI��<.C�$�~��Թ�d���}c�5�-�QrKKMF�B���+�&?��G�6SJ�,T���V>�Oy	Jھ�R�T���6�_��}�������ˡ�Z�gt����Y4� ��GNg�ŏ%�[Wue����nN/���Y`��"�-����v3���mE�lцQ5����T��#M�-�d}���Am�d��@���
��(�N*��DF*���NU�+��&#�P�7 x�4��o��&���fQO�g5�.S'��H\/>Z��� ����+��-�+�ג����(<���l!��(�p�%�C�H;}��hΦZ86�C쟨�՞h�+nJZ*7w��k�(9�u�Nȩ�����l>����h��������9Bw4!�����z=�w��kI�.>'5�JnՐJ~�+ĭ���6^��n�����U���`Ħ%_4;�N}s�A���4��O�%����!�Ѵ�~�|��I��q�h�)J}ۇ���
����tT����+��M��}!a-ƐòlkPq|��Qb�N�bn#3c7]�����"2H�_(]��Hd���H(�́�xy0�C����;���'��x�2�*����	���.�����	��'�3�M�E�Py��_�=��M���7ײ���#`|(�$0{�D��uR՛�Hk��l�.L�0�H���)�4��뚓�{���Q@�`���YZ_������2�O�G!�H���$�n�y:��A"(��H����p�����O9��P~��?�-oàS�X{ ���7%M�=Y�W�dIףּkjGN�\P�T�<d�^��E` ��y'T�ݍ�3d�U�d0W�A��W�'�h{��_�\Cw��v#/�;���pn�V��#�EbBk|(^OY�����b����w/�"g嫳."��kN.�#�͍\J.��r���y��B;TY�Ir�H��Π}�y���l2�10,,�p:'�)�TM��-�t�h�N�"�*��7��"��u-�@?UJkucCZC�ȇS�N�76�>�I���k
V�S�.�t�8��P��p�W�^��,��%'ګ	��>�M��l++̘��xm�BK��q<Ra��X��
�.�v��i�p�/m�lx�Y
��y��7��f���-����0q�=z�Z��ܾ!y�'�T�T1��C�&��iR4РNp`����	p����=oB��d�P����+N��J+�t���?�k�Gm�[U��L	2g-�	|t*d�/_��ޥ�@YSH��e�k�������a�.�Â����h�ק���VRH�r�1I�\c�lw�Q�ۇ�0�,�����V>,u��~S�zZ�8���/�����* W!��}_���՝ѩfy�b���`��ⶺbo$�dNΦ�|�"x�J�:f+�@�Koq�_���^tl�de���M�(��d�9�%8�j���� P�$_�IN��*���BFb�cn(�-��6�Z�.�w��X�+�?Ce�Wωȹj��f*�^���o���6c�䝐Y����r�tE�R ��1���-��ॗ౱�:ۥ:r���\�L#�Me! *�	v��_>O��ES�W]ھa��
�9�&�(�K�\5���_p^��&��+\�ҫ�s��X_��b����2�>���lM��.��3!�_c�!�Rh�yPXEQ�o�J9� ��8���^Ts������ɂc�مD�0���&_�ZG$�
�
��j�*z��>��hp�>#��T�ljiw�J����âX�s)$a	����;io�|��I0Y{���A������ ��?T�� �@;	I�@���v޺�}��/�UΜS�5H{��7]���>
	6"��|a�
�6Ɖ��������D���oQ�Y��	�qG�(۾�z��r6NaNj�X*������WL�gc	��)c�G�}���[MKv"���R������1�Ъ�􉛺�!���`����)�Y��WʖPBC�9gm��2�E��#��`�X�fI4��9��1��(���F]��>;p'S��.�
>���M��� "�V�sd�۠���!������y���H�i�3��a�'�����;�n5ݍE��Ժ-s �W':�q�?�0�^_Me�Il��"2�%ֱ�vt��0 �Z����ܡѹ:7��?�KJ _�?�˶���D��#@���X
C��(M�3Ӳ���
�LS�P'�������2�*�q��ߜ`G��eq�|������g�w�Wv��|���������}6�@�v�Q����@����(��F��J��h$Ėw󣮼xA;�/�4�g#b��G5ވ��~p��Ak
�xɱ#d�l0�'�r�1���R��� e��LJ`}j#���3B����@Siw�8�F���A4�<H������<O�e�1�([%�r�0�Ŝ��t_�����w��I��7k5i��zG��-'�L�aH<���c�lb��❷�m�-/��X�
�Hi�f&�Hk��3G��5x��S�����E`ҥ`=�Zf�(�_f�qP�t�h�������N�N~��c/m=���R���f�WD��O��aⲨ�N`SD��T�'����C'd�KDg��XS��DMM�����b�^�d�j���/��q�{�qS�zX��M��L�����0�9W:������ E3-��^K��0�ۇP:E�-FO�=�lPᑳM�V�BC�l�bRO܀j�Z��?���t֟���!/J1�L�9+�5f/1�0Qi�7�%i�/ͿrOg͙��D�_�����A�o�CH,߾�Igy��W���(�]��G?Q�����{�M��*���wyaX^G�	�f�k�q���b��AG�_��5��'q�3>��ѫ����ϲM2�����y|�Ȓ3|�H���[�ٗ}1���y�N	��M�Ữ}�LrJcJ?7<c+Q�NR���-\t�%Fp��kqZ���J��'Z�ʬr�v�~DMꙮޮ��V���#�o��#�|h�S$��)Mh�⹆��iH�6�E%����N^�1�j!Q�~>��e ��e����)W�6T��)*'A�"n36H��&"�A�٢:�v�d�"7���)��;�<�ѝ3_I
JE{�3�ʂN:#�<EmE���8_=	q���F�J�2���_-q�"b4�J�&2�	)S�:��041�S��eV�C]<�����	A�1R8Ā[ᮖ�Y'!9�apv��)���z��K����a��wP�Z�dt�Q-�R�(OC\,��F�|X���?6]�QvU1IK>��.g�F�$dm��_�<6O���kP�Q�����Ҷ�v7"_�]x�G~�~\T�b��\��]�6d��P���N�\���,I�}tR��Q.����-��@���z|Bў�=x��j��̂:A�痢���V�da���g�5 &�	�]����9����'�Q![�	ݐJ�%ȶ�x��&s���������@#K�j�}��u�.��r�q�4�C��yza��<I/a?V��Ou�{����AWW�NL��t�S*!�'�-��mLG�>_�&��a��Z�]q�s���`�E���q�f�~�HF������Ec�����~���0SN$�%��XW�_�U&0��0����^8gR�Nf2���ԗ�90���a0�K\�󉑗�%_3�xvۼW�;�� ����p;���EV�}�E�׼i�2��Zv!kA��Pb��G�����Î��^�E���N�?tf�QW�z㮪T�C��RUOPuk;�v�)��م���rے%x������Ī�zfW���KZ��-�y�o9��T#���V��ھe�\ҟ�	l�M���b�L��s�N�<��|ݵ15A�o��k�ט��

]?la����(d��V3Z�����T煂�&�e[��V����5�q�,˼�^�����&��h�-���zõ�b<���kkH�ӗn�ث��zl���`}K�e����R2+���b78�Z۰�bqi�ל{�I~��'Fu�Oկ�_�2�)��ˆ)f �\s鐕\�<�g�:{@�kM�SW��^s���m*���'�Uw9B7��	~$]Dc�C���51�!�Bv�^�8Hz�����4MS�?�~���1�,�o��,i�۶�<LX�Y	~fa���u���2N{��Ö���(=sc��Ą��6�eE�!�n.|��H�y�����&�a�f���� s�9&E�3i�m+���z�UEҨ^�����(���3�(ak�K'�Pܲ��J\a��3҈ 8�!�M8T^�W�u�y�'ޅX����
�.��z�2p�{�xV�b�?X#YK�FP����7,�lx8H �k�j��#*V�m���.2���c�L�b�:�]Ϛ�h�<=��
���ͤu��x.����_�rh�"D��.�CWFF�l@�m7��q
��藛u��no���B�=њ��U?|�;]a8�[�w�*��\�HkLR��
���H��w�RU6�ȗ֍�)0�>�
���{y�ܰ�4�&���a�p!Cg��Ј�0�t삝��)�2���y�(Q��>���b��i��-�1����B�d΁.)f#���,ި^Q�k>dJ�k�S���yJ����<���s�	�m��/�
�ŝs��UJ"�+���V�(	 &���c������ Z0)Յ���V��_�P|J�/I�D��J�ڸ�FL&'°,^Z������g
On7�+6��K�Z!ϙ�*'ĆR@��+3�?r�wy����^�8`�R:u�Vz&�@.�1y���Z�:�p(�Ȥ�r�_�/z۰|	[�jNN�-l�F�i����[�wW�x�j�*�m��B�b	�*n��&�
¿�`��}c��-����!̎�� ӽ1�c�@�ߨ�5{xj\�l)>M8�.���_|XHj�~-z���0���<��/VM�r�(oi�����²V}�g=zJ�.�ra1E�]�*�s�
�i��-�gj�suZ��/q�U�괛����F�Dǥ���<Jq���x����ܐ�-&<���쌭r4}td�4�>2��M�NC�;���`�>��V/��Q$y��85��~����F�aD�S���/�oṤ���7ѥ`|Z!I5;�t�k��,&��BIC�Ў&���P���I�*�p��S�+�*͜B�P��N�=��� �������S�����(��	{��~����b��W@X�؆aBt(F����v�*�����3 ys�4�M<G�Vx�Ⱥ
�;�c^0;5��pۚ {1����}�Pnrw�U��	�^�i��:�1�WU��x�)�Ih~������r��Ɩ��V�#7���LNV����`�-�Y�DGj5 ���57�ܷ�nܙF���Aǔ�=�������3O�Gazo`��r��o����&1&(�	��݊�2S[�E3>��!$V��֭R\����xe@7��ys��H`���v����68]�;Ø��)�&�'���,�b�rX�0�0��7�kѹ�o��l�HZ�˕-���D�F�O"������x	�K���,�%y���P3��`�_��ޜ~AoU��e�V����ߩk�]`Ca�t�UC���&�k�%fj$;�{����u�9m��5���o1�
��^`˺ ��!��H<�6Z��9�H���̪DA�Im��9(�7좀Jaοۙ/H-h�&���:s��AT��"&�Х�}�q�$�������gJkv)�3n��pR~��ӌߟIa$��㻭Bk!l/{����zԝ&��o���h>0�S����o����0t��>�#�4od83�N�P,�a�����	�S��{b�~x`�C(0ru�;����Ӭ,3s#Yu�CTd���S�?�$�e�pb��a�:�	`����6� �BTy?T�k,͆U����/���~iXlxVHYEB    fa00    10e0�p��C;��}�<�z�ޭ��W�M,d����I����QL��h�GS�#0 lN%�5!����/���3^��?,�鯍�*ߠzo�l.'/`��Ԅ�!Hb�F���s��1�E�~��B@2����c��{t^�����׭n�u<���y�2uB�~�>\�!�	}�#��o=�E>���돧���:��_O8��� 謐��4��d����$aM=7�M��B#)w��v@(��c�?3!�\�w��1��x�]IBO)
n�@yi��~x�`Jq�?MP\���6����#��a`&����3�(��u�~OR����K����F?x���Pv?6��� �}����cK��X��^䂒2�B����S\�%сW'��b�EK}%�ų�7�%����'� �"�p�B.�O1 �i�		��u\� ō��fQ?B�w}���.̧dC�a�$��R$oS;�WH3?M΁��|�A�o�]�IuӴ�-B�0���z/>�G���j���M
:��H#bX6�	/�ja������ܞ�M/��̵�dW������z�ܓ����ipij���@���gen�6��b�uɡ���^�)5������L���������{��u�v�����(?6�%*E�����pr��[J�Ë��8��o��QK�-`d��}o{�����p&S+p�s']� ����{P�erѼ,�>�����^KYqPZ�������9wy�aC��Q�����ڢ{/���Mċ���g�E���O���.:��W����'����[C�2��t[j����+���ֺ=�\��UkO��)�f�u7�7gI�I���Hg���pe�>�YG�T�(�@IwQ�%H4=����RP��p����)�0s����5��:x�~=�M�Z5�$��C!<��m�,��n�:
� �srv�qE�INf�9x��z�I����c�RB�*!�q�'�Rc���[w�.���s���jR`�I	�:m�@�-�L�w�Sq0�kWv�YQV�y�0�I�פ��_��ྞɌf<��k��=SK4�G
@�4�&E	�����es�2��5T�8fb·ohf�I/�u�T$-)$�w �s�����1Ώt;z2�xﱶs��d��2!��1a�C���$B� �Ƃ{�sF��f�o�G:Om��<��M;-�~Tb��^!��c���V�ڲ0�IYf?�u��x��
�Ғ�7���9���J����7�Ǒ��Y72���O�ػ��P�M��=�4��#�1*��F�����X�`7���QdXh[q?�"^�@�"��&�����[���z�9_/|�\���� ��%��k7�_	��;����;.�1� `��V��Y�I���4����}�|�'��h��}>Z1��9g6z�����QN�ݿ�x���f����#�L	jd�-����Y�>�"G dt�4��v���o�#��]�o�I���6�������)�¦���)3����f�f_h)*�L��n
u�:�	�)&��׌��#������rٿ$��t^��Mv8eV��R|��=*�u��f�ėx��TL�0E?�e��&�R벛'h�S�����^v�J_9�R�N<ş��b��MW|����r u���WMn�p��(��ؙu1�Ń����)�8iq��\��#$N�O��.��(���`�x���IB%�&|0�e1���s�
}Ĺ/xQ�j)D����Dp�N�B�]}q+ȂDd;��s��,01-�=T�h�=��[�Ņ����EԧűK���-��5N㙃�����sB3�lQS剑�FY�x�0�v�M�K�qu���P��t��B����f�[Yn1��D�e�daB��ApY-9G�����Twk��:��ǹ�Q�`) �!'��M�|���_��D�O�����N��
�e-*2N��L���Z;4M��d����ݬ{��UL�3�iH�,�h�Bx������J�0n�g�����M� �lxomo���t|�6��v��s��^ĩƓ]�Zr��r�m��D�ks�H��a+�x�)@��m��Bq���W����^���N�϶i����*1�c��-�L��&�y޽���Wq�B�
�P�=�h����>h!��u% �����y`i'q*�嶳o���B��O@����Δ���0V��6�Ⳃ���?��/"�<�P�A�a�&�s��'�m��2(��'�
ʸ%?�1dX�W�
��x���8|����s19���_ �@��;F
\qX���X�������)����TY f�i�,��@�"y�R$&����������&{W.Sf�,�>u��Py�S�Ɗ��g��A���!�������f�8����ّ��rk3�������{�JI��l$
!{��+��"�e���E}�y��0���Q0���,���V4�;ӛ[j���>��𦶹~3�f���e���o���cP�\j
;ץ��+���ϴc1f���˚!a.��ٷyJ��r��y,��fJ�φ���$�<��"��Ÿ�C�J��!=�]_�@���s��AvI�"s�>�O+��#�?�/!gL\�0�X��~X�k�!�6?D�yrc�~]$D� �nMX��5S�_�E��X;�ϿL�we�~�)�-H�����?L�e�m��</����)h'BEA�K e�.V��z���^WbcS�h�`P6�V�f�!e��Fa��s�`��Y�s�ap
��
�_S�.x�+�b��Fu�'�� �k
�x
z����3�ޅy����d��DI�&�ҺY�,�_���x)*\6MRQS9,c�>����L�I� oy�#���,x�5�q�U�g�
c�F\�z8P�����0�5+&���%�0�:7>S#��[�r5~��:أ�l;l���J���L>+�Sy��
��}���� \���c�I��eb�r}����G<�ȬqQvǅ��F��UJk��=�_�����WS�TYހ<�90-;���[��K�h�'7��xc�۫#��3n0Ki������!f1��1YT@����_�>;����))�Č�':A�j�g��M�	�d+�A{)��(�BU�(X|�Bp�?�cgB	2�sR���6��&ZK}��p�M`�r��U&�g!�so7���u2<��0���ŵw��&��R<M�Z��9�|đ\:���7_��$J�f�wC�5��E�O��.\({KH�OOe�x\��/ȼ_���ڢ6E/��e����!�P�l~c�g�'�>5>S;-J�����	��7���ڛ�ʛ54��5�e����VݹԦq�)� Zi.�B;z�9��֒��,M���)���9�y*pM�f��P*]8�2{.q�&Nt֖4i���k27����F������T*� P~��4˛��/��sOR��]��e�>�{))ON�h1����N}/�gb���0���������U.��Vc�����}[�����Q�K<��������h�'y$���:��<L-�3;��@q�}ɭ�Fz�gu ��_/��q��.r�%�k0eU�!��B ��CJ[��0��Q	�ꖾrtguVf�A8����W���Ă{�r�@�l_$��*�5.Y�/�ziu�R�)��ێ�-��T�k2���5��_V���v'�I�*�|��JV�n��2E �e�fH���͎���=�S��=�W��&�e|�l<�Ƃ�q�9 �x{b}�b���D:�j��X"�!�֒V�7��,�$Ҝ��%}>�mk2D�nє��66�%�+}d�q�w� �g���ex�.Ą]&#L�H�e|��Q�b���7�6�k@��:I^��{k?O�eO{5�*~�O{k�$E�%_h9�cn�p'��i����0h�-��� d����z�Y_z9�U�� �i�گ��ľ���o}	>�#"��<�gK���q��uŐ�4��ԋ������V�x"�����ϿB>�`��:��Sz!Gr��i��56�a|�Ή������u�����V�Ĕ;`	�R��Kh��m�������_:�C� 0��������)�l��@�w���w�T�,�rƌi�̽�U@��1ڏ�v��#�}������Z��@n��mB,�܂�	]�º�Ch��q}l{p��M!�'��w���6S5��s�}5ǌq�%J>Q8Hһ.�F�F�S0���b��T����z�(8��ţ������̓�H��K�U�`�-⡶,{r����fo���h�09�XlxVHYEB    fa00    1860N��:hy$����.�GǍU6����>j��23������p��-֔nm�$�oGeUi���|v.����Π�$s���mi�'İ�w-1S��jȑ��O>�I����ukS�iC��?�x������@Ѵ�IyZ�M���(͵x�f�������?��H(��������r���
%�?ɥ�U.�᥅~jac1�W���Tn-�?��u��-r���t݉�"�vZv�Y�[Q9d������Ȁb��0@�}.� G�jH2T0�c�2Ǹ;|�®��,z������F���Rl?��_ ^���Yx2�o�?��z1n�����׆ƹ*��iۀj���8U�`<��'!DQ~5Wԧ)��\1��%H*�o�o�2fn������1	Q�ȿĢ���ˠ��F�j��=C璇�oi���1�eudg�d�!Y��b��/�A�.vX�iVJ�di�f��L!�Bt^h5��U�J�MlӬ˟��ܥ�x��gksغ�R9��W��r=u̫���| ��]ގ���Y���Q���ע��du�2оi��l�Z�M:9��>-����d��׃x@�C؇��*��Ӊc�]����ϲ*Fr�Fw	R��̮��a���,Qt>��e�������֝ћ�i����r��Ib`s��-�3B�"��+	Q�(ָ��D6P��xո&���{[:-Z�/o,�e�I�
)�C4cH�d�t�@����Y�	�d�Q{q`�@�:�CHl����;	QZ���FBt�#��o����x�Q�D��@1�F�	~�z��;I`FvM2�L�4sv��i�� �l(�:j�Z���ҫ���wIܛX��a��*W����\����+�\�n�p�yA�}��lE�6N�4�U�zB<�v+�]7�¨S|-L �C�Q�G龪	�?u%J�}��<��L�WW�Ɏ�9䋾}��@���߻ҩ��#1�v}u�[�L�K���U�T���w��Ƞ��Fe��s< ��×|;���]�P_��	x�W��d͞�z�v�����'u��Xۇ� 8�t�7S��-s����Q��hD�|ʽb@�('�$��tK���q������O�9��F��zd)��o���HX���ӻ�5���B>�b�t~��{��O;m�>3�Ui���~��tH��M��"��!�����)�����mh�5[7a�,
�o�e��X'�aer/�s���	kĹ��7�p�qAz�5\S�����8l�(q�D�d=��>o�j�9s"��h�i1;�'ci&m�b ���
�����rL!=Y(Zf~�a���?H������&�Ң� �6߮��o.	����핊CVy�E	k���4����z��db�T�},�s����wy6{��F<{�!� �O��|F _\��y�0?~g���.3���QR��o�F��4�/E���%F*r)+��A*�?-�E���K(sW�I:<u��C�#�w>��Z��/���6p�M�2���#W�(?#���='s�#�Vܫ5.��#w�	���n�	��T�mC�C�i���ퟖ0�g�ՆZY2-[=��/�����ϑJx��ش��c7l�6���eF�ӕ����� �`	��gC�"�x�k���qx��`.�
�Q���dvr�Y0���/c&<�r�1_'�n,.�"��:o�y\�xS����.��p_�Q��X&��m#`�u��Uȇ�H��d�:޳G��	�F�pul9,5��Lc]�K��$�5�Y�ٹ ����� .�.��BJ��N
TW���7iB!��ŷ,u�ݚ��%�i:�Ba�V�t��v�Ӵ'��z�h�mB�ĕ�)�]c�@W�ds@j��waO �x����
�@B����l���0MIy���GO�{�U��Г��:�9�xײ�߿�e$�k]����E��w..y8f��핫6�����V�7V�"��v{��98�9�S`ST�M�?<����a�+�Msw�=�9i�m˖����h�8�&s���%' ����J}���	������[�mFەe���H�\���=�3���Ŵ�ӹ猅�A`�O����dU/�p��b�K~KD�&_X�2���W��9�x�����kh#�?���B��+	L�M���i���I��3l�9�vŎ�^U�p�e���.6)af�f�PqRC;�@����?���������-��K��)�=�[��/8B��fj�x�L��s����L��-Ko�ak�&5��p*��4��n�I7g!����"���xę (@�o/)0	�"r|sݞ[���w�����p񟌍�lxnЍܞv ��K��\Y�_~��J?��t��-�:|e�I�Ӊ�m��>$4�9�E�ұѾs6�š�Xe��z�uj�!�H����5�rPC�%ؐ�%�h�����MW3�3[��+������x��/�r#m�� �	J��xX��e��������\��&�5�0����0
��7���US7H���˲?1p����3f�y3?C=F
�#�#q:�Y���x���[~g��|+��ja�I�#�?�=<�4S�s!�з������R��B�kjR95 �0ޯ�9JC�� Q�#D�y������Uv֨���Ⱦ��9�kXT��z2!60
�L�C��эd�I\�m�ʸ��[&�s<���Ȑx�s�, �ш|&�E��z?k��8�#��خl���)U{��ВAuXY�Wt*�ǝ��z�d�%(#�aU�O\�9�*)q��r��pG1DC!JL�X9�[�0��F�]��-]d�^���T� ��ֽ�)���R�H�S��f�p��|�g=:]8|f������a�Z��9/�H5a@��c)�6e��u������>P�Xm�A��q���5���)��k�28/���f���-&�m�ƇvMhR��;ȇ��+�3l\O�5s��P�SR�Cɟ�0��Ϋz�:s����?���dĈ{���LY|Y�)��-�Ɏz�
}�y�^zR�;���-���3V�5cSț<�A�I��bk�C)����T^k�hs ~���w.�qa��S∻�~�> ����L�Y�*g��c���bd榆T�+|�ϗDy05�r`x�(�O��~c�U�Q�6*�m�b��S�U����x���I��a7�h�Ty�E�=	P�Xcg���[�K.HJjLy[:}<W��f+k��ð�q.�mh����M,��1s�/m�W���DZ�:��Ѣ��҄%+�y�Q�jMq��M�����l�-du�����N�_���o�Pg��S,5^�t�Y�Ȧ(C,d�6��r:j~���i"Cޘ`q����|?w����!�-]�w%3s�Qf�$f�������X���-��5�j7Z7�^~�U�$>5�C�pM�^g�p�u�&#���H���~%��)�d	��z:�%6����+RJ�4��<�c�W�Nʐ#�j�E�?�F�,B�=0å"dʊPTn��q"�!d��RMa� y;Gfl"�È��&5Qr��k���=���}���'ɜ%T���^C�h�Ѩ�b�N5��HaW�(��崣&&�܂J���@��� \�Z���)�8	
=��,Ө���#�N�4eܻ�)�:M5؁���I�x�z�m3A�̵)��8r�J�?ʦ�%e�w�R9�=n�!^>�`(D`�5̰�)��
��J�2�@R�{��wax�Ȝuh�*Pb�h5_���e�������B�O@�m���ϑ�̰�^L��=����=��<���Q �9F�U�e���g�v���Q6�� i�ޤ_��1s��?~yv�6x�*�q�AV�#v.�>���XT����cJ����RY��/<�K�x0q��}	~�pyiA�~�\��c�쳺�ر�ۡ�U��_}R��מ����0]U�\oc�l�q��?,u����@�a�l�x�z�.�j�ɺ��BwM�Ϻܗ+	�R�S�`��D��~�H���>�.����ǂ��K+-(S��)'y�<�_���u�	��*0�f�)�Ae�^�lK�j��. �86������$$��eG�ዿ?� �Ħ�;�!�$D���A����}��7�����r�V��rVp7���Wp��ƷE�%�k&���f�R��Ͽ`l#����9��	9 ��w{��jJ�F�ș��+����:�p�FG�N�s��R��_� �'�\�/1w5".�"u"d��AC��8�+�b"��t8a�����'�>�s���4J�:+�����a�}p'^e�V�V̶K$�@g�=a֍�zO��>�"�@�TB���b�[����{��:��C��c���8a�AZ�ocNH2���y�-�^k�ŉ��{w%EV�v2^w���Z��	�⃡���B�F�K�AK��uq�z!xSiɰݍL/�><�ɴLl�����C(��N>�?�ȉ�r�EڟR�7\&ѡnmc��g���bv���6�}��w�����%�}m��Hwˣp�VO�y��k�?��a�_���D�$6ku�a"��¨�񆄅�~�1-L=G�L2�����ԉ�����Ҩ�ϥ���Tѝ$N�j�9�ۘ���КZc�.�}����@�s:d����hw)q)�e߁�3�����|̵�,��goB ����L�]6L�זɹ�@�w&~/L���-��VEF���0��n8k;��ʔ��'�Lͻ	��m���Pp[T�SwO$��i_p|���2b>�k|�M�H�P	�Uc�*��h��!U��L)��Q�/Vl�W �R����5״˺��ddEj��������� ���p�=jj�"KL�M�U��ZԬr�*�A�aAؓKa$y��l�i�P��X�s^�*sUu�W{z�$���%��߮��MHa�EE��,'�>y�g�/~rY+w~���3��ˇ���s��C9�-_�٭Ӕ��q[������EAAP���TW>�9V{$U�����p!��r(y߄����x�6�ۊks轂���U�~��<G�>cs�;�?��3)֠��U���'}N�ƕP��7p� t#���C�r��bN8���J�����5rR
W׉7�M&k��#��XUOv�	Ϸ��2��='�V�_bF����z���ʮ��q%��q-@��B���٢Sa�>G?x�IV�6�����=�l���� �D�D���������
Ej y�Е�r�/'P���oB	���N�T!�:Hj�|������	ܲ��F�����Z*�=�(�������x��Ԗ����å4�wu�EL��C<����P�LdN�Vw7�D����W��L%{�I������&��4c�7Y�G1$: j]A���Pb;�/��0���@e��q��o'I�:�E��+5I'����6��SY���~W�8Օi�kEq�j]������F���􀿧Ľ�U��牷�:��z}&1�f��l�l���.�n=Q�����g���zl�����I�D�se �e! 	T�
�x�����_b� ��Ӑַ;�i3e�=�������?���X���!\�g�z�J�@%�XC=?������!�/\���Ț��7���L�q��V� Ϋ�� Pz����\˄H�'J��r+�|FS��ӻ��99�1+7�0)��F�g���T6��l^p�Xf3��G$;Pt�����Ȣ�ұ����H��m$K�0��l�~siנ�վ-��u(s�1@x���Vƪ�@u�M�`�������-�M��<3GDu���Ѫz�ߞ6��]l� �jT�k*�~1QS��s�J0qM�7���a|XY���s�Fw2�������Èk�8�;�k|?mN1���Oq@{��"�2!�,|���9�����4S�� $��ܐ]�����N�-;�Z������D�Ֆ����]�܈�]T�����Z�t;N׃� ��A	$x����LJ7�R�����L�$qts�>����/��� Q���.�@�8"��ڝ�/gM�ϼ��+��U·g�T��ijW[v�蘞�l�-�(s�i)yMS�-�$�5}��Ӆ�ֻ�U�2�ʺ���ʯz��P�R4��4ueat�K~�'���|��02��ZU#����B��{w�v�X��[at�&�3��P�"�!;�$?؏v�HRc8�W���<H�dC�<���
b,o�9VWE�8Kc�D�[�u���VXlxVHYEB    fa00    1720�N�v��|��崪R̂��� ^�yf��~H}�K��" �3֋2�gm�0I�Φ��=�/ٹ,ć�h�VD��T@������p��	wP�d�V��������3���@t��EX�jc4���	+0�Zҭ��7�����SHu����,�3�VD���ӟda�E����O]������GҼ��V�V��H�^a���bE��u�!$�_}$�7�g*���fXȪ����<���,�����y�a�W�<t/������Rα���g峐-b^+9=�j"�o�7�D�G�����ɲ���pg�	75�h��'T�����t����^
���\Pk!������nf�//����d�!d�!��Z7MX���ĭ�Ze�Ț��^���h9�� 6z��� T���h7DM\���+ET���LE7-������Jj.&yļaB߃<�V�������#Y������'���+خ��/Ty^��1=K�4gj5�jP�]Xow�!���@ZH�w�x�"���d<�x���z_r��O;��v&Ef�"�n�W�Z�\ی�G�ߡ��;` �h�l��"OD[H^�h�ͼ�&�PL�Y�I s��?Ww}�
z�<lQ��-�MG	�����Ps>*�m\1�\�,�㲶�6�/��!W� �^}��>����$ۧ����������Mu|��v����X����B�E�fc��N{Nd�e�Kކ�Sͺ�1��M!�
��Oʴ,*z0�f+�c�u��鼂��k�ky�`�it�����(�P�{���9���?�d5�����G?�)(�+A��X�̈́��<f����_�e�k���e���>X��R@ک���������G͉"A�,{{؜��![PP�9XC��zZ���r��bm;fu��Y6���o0rQG��?.�89�����:��St'R<��`����☡z�gJ9�A���7�s�>���l"FmҼ����X��#[Y�9�`yaP��k
�U�4�Ťgĵ�*�,"'P`m���ў�Wb�9��]E� ��P ���=���=����Xld;�ɒx��<'��/�=)f�^�Z*�Pv�y��hǖ�N�DL?�V7�E�1��S[�qa���#Ώ��E�n>6��z�@�3��bYR�Y����0Y�[̡߭BT\(��3Ѷ�Pwr�k�Ko���ހ��vp�)��SU��9�=l+k7���*ʡ����}}�*�uj
 D���{��G�&�H�W��̼6���;���F��A��gL�=}�Kq���������+�,��l��CG��(AA���M��z{��f]�ӏ�����|C:5$5�:jVn?,r�gc��e�F���B��4���+��X�
;�s.G������E9���Hp+e��*:ǃ���p٫��-6��[Rc3w����XY���9��O���R�,K�� �Y��3�T��U�[�G�#>W@��/�M_����_"������:岸��E��ʼ�S�}b�9�ClKk={gu�-�FD�+L%�
5���'�P�c����=ľ+kE%EIS�y8q5ޢ4����j�>v:��퓾�q����2�q��a��@$.��Z� Z���i�NO��ȷ�6AZ����i ��>��%s�.g{hwH�X���w��I!�HI
r��9	 ����s�h!Cb��ׁ$��`z���*\֠��eӦiX�;�r3�u��ݪ���+6>��$��6)�fӘo��l��T��ń�sk�Y���
�|7첶R#Rd��Ý��TcA��K�ΏGu�2 j�VQL'0�M6C7��З�Τg�Tg/�1�Sqq�r�����~N�m�&�
%Ƥ�&գ:��O�@�]T��>&	/p���"���vzl�U�z\M�Kf�jVgN��\��v��T��1���>���?U���c��1�D� r��U �g,����CP+��x�,�5�`��۶��_X�7VF��Vg�ק1�w-��M��A7���)fg�@����M�oW��I6�����Q�g��Tŉ.���;����.9�2�KHq���<��4�MЯ!��4���vO����U4�_�5�?�`���a��T�w�Df���[�5��K0��� �L�oۂ,�s/8"�T�].@ r���XU����1���ĕ�J�2���g�:����t������W���sZ)Z��,�h�����I�{z���4,���x�W�ү��gep���
�/H��k�-%��c����H�j(V��3P�� ��x�[;o	�-:*��y��$�k�o��2���v;��@3L�	�bʋ�]���
�It1�;YR�|7J��|f���,�K�txǫb�(�F�@G��$���F�bg�B�2��3+*$�Ýb�P!�6���U�!1JL�q�=�{t�;h����P��Ǹ��`8]n�^�^�I��qn���}}p���6�	Zq~!��Y(�|Wɢ�����M���QU\�|����3�U�x��Z�L,/'���L���ϴw��G�ȟ�y���P ��x��ىYw�4ٿ漑Ӆ�j�Í��͌;��B}�;)[��e��,��y��l��<(������9�AԵ!�#b`	8!�صLS@�/zx9gJ7 �O��3)��,ig
���,4��2�?Z�V��U�杻�f��[yt9'�=e��zŬ,��;雋=�̍�'r,�ڜ��T��?�ʬ ���2�$�з���S��$����8 �e�h�>��#��*jW�3�K�O�|^PwS�^'B*�����J�Q6�kd�o6�a�Z��Փ�v84�.[V%wΓ�~8�(�]�A}W)t����j�څ��A��m|Z�f�������K\�g�)A�D��M������Q/ݚ��V�tJ�\Y�>Lj��\-��E��|�;ĿB��fY
�BEdu���D�D���O.�B!0咶kM��\���lԛT/��������4�"�f+˔z���������Qɑ��Q�C	����I�<��l�j>oy/νvN�:����NO�S|lM�V�j�ǌ3��qO��pm�E�Y�'�_�k	�&bTbqY4f/5� �G0�i,�a`�����!6�vjv.Q>u_�⫷���-o�v|+��-j��~gg���yB�4D�������P�{si����S(l��A���D���3#�`�GkX4�cj���3�˯�o^G���w����$�©o-����T�_�)p�RN����"�%#��p��	]�ET���R��wV���)8+D�¶��lZ��#���v�)f�!��<�둎�8KW�J(a�$铫�	d�����@uL/WȎ����A(���!���K��Z�˓R��e]�y�ߌʯ��'*���l��
T֑�Q^T���ǹ1�����3⛗�"��_Q,�M��%U�#��nUEt.��`Ԍ��mVE<���; �J<��o7�dd�K��{�L��K#o�]�r�{P��wF�g�3�VY�`�����P�K}�t�(�!���}!�}���WB���94&&a��`4k��ӑs��(���ֳ~�I-���h,$(��H�t&M�S��n2�ձ���^���!3������#���Q�X�G4.����!�����2;�6���$L
i9 ������ ������PJ���G?�u������Cx#���jS�ޞP��6��IPn�2�u/���A�9�nFn���6��	.I:XKm���@<����'ĸ���,�N�H9.%����M1�X��`�ɸ�d���$�(��pM�3q�����!�m��Z�pʾ�0� ѥ8L�w��4���`u
"J�ɸ䢝�]���Lc΄��>l�y����Ar�|��� �es��$Ź<�:Ղ�D�܅� D��Ŏ|91��Дv�A�]��Ԗ[b,�ekq�
��y�\P�{�Oi�*xn����s���PP�}�*���I�g�|_��1�f��Ũ���#GY�]��M?������F!�?�eD;�W��4&:BW��x��U�u�
��|�c����,;&z 0�>�(�Zs�Ҵ�jQ��������W�&Dh�kj�q�zu�5��(���}FX�SjG��� ^�jsFH�x�}�b}�gm}�J6��S'6�F1s�*�K-�T�,��;ʕ�S�B��^���%�a�˾d�ڐ�4�xBa�'�r:�}���l���ߴ�t��h-��(����'i{��M�4�3m�i �(�Y1y혍��0�xكf�u���D�����]��2�WK��^2�-ʄͩՋ0�<pm�O��2y��~���^/�A�Z�vE�9`�M�
k����S,�*i�{�3�	�a����m��TM�Zq�&�����O�_̽�5��Iv:nF֘.�94k��8�d-Tf��޾�D�2�����T�lu������?"\bէ*�@��y��k�|ē�a�T'r����;+B� ̯�L/�:�䌮!��Ė&!Gڝ3h��[!~hW~�|+3�P⑾�z��Q2�)������a*�ݢ;49�cwR��#�0x���3ݫ�2mѣ�_���.x�jn��*�R=8�]I�����u(��N��]����pgU�E�
4��%%}鹘Uf��n/��ZW�`��C;f0�J�l(>�,Ҙ�(P������u$F���%�gE��ȯ�I���^FnP��ߡ�j�U���zb}ղQ�e1��Y�s�s1����?D�%j����3"�������ѽ}-�n�/�1PZlF�u�d�"�n�u��xv�Ʌk���-O�N�݁�K]vu|8���@v�(3_�WW�(�=�
�-P�aR�CD'?(�e�p�(v	�הi��|� "+c%A�T7�������:��I��!�BsI��*E`��+4ډ��MC�_�e�<pD������C��K��;�����8,��U���j~}2�K�����"/f0��`0ϕ��3-�
0��t�ҕ�ms�R�P�:���0eCÎ7���9��c�&���cvM��0س��N{|���f���T3�Q��rbL����ƥ�P{�-彴)gQ������4���ׂ"w�'MDn�i	�90n3�~�98O�W�;KV=""��6�!k���,a�}��oE��<�_wq�'5�Sڄ-����W�D���d���6���W��ʐ��^#y��n���C.��6�)�N����{]N;��/KKcSA]y#<��՟3���ׄ�XT�4G���Lǘ+�dY�9gmN�A�0��8���WE�k�.=�t��I9�
Z�����n�:7��w`]�����F��`�$��*�	߃-�K��5�0�M��
ɋ�~�k�0�+��=vT�/�$���3��L���;��*ݶ*��5��q�P7P���0)���J)	P�3R���kȿ��R\�?3V��좨zڰ4��Of�o�,4ה��?��v�E#�.�]�Hx1��Bvޜ���AP�W 5u%��j��ۡ<�i*�V�Bq�ʮ�A�
��Q�4��s�ZS3ˋ���$K�u9��;3�q=Ԭ���y9��**���ɾ������`و�i4y���gw�~b�'�@�ȆW�<L��a�4��61���LŌ�|5̂��!'�8���S>+�|�D��n��ח��M @��^E�FY]�8�俉7�'��̳�T���%�'�c����(�IJ�A*x6C�X������˄�[�G��~Jw{<��Y�'���ؚ�D�V���∑=L���`��K.a�6�R��XlxVHYEB    fa00    1500R�D�٤��$y��'"��c^E�{q�W�u��\Gj��lᰚ�C�RD����"p���q��GW,�b�`���#4-H��u����Tz`�0�Hv+���Wm�^4�x։3��؆�����ndq|�,k0[�ԟ|��P���w&3�x�F/�^�
K�O~I*6�4���.}j�hX9;/qp�׋(M��lҹh;���8K�z%�m��
@j�N�����&�� ~�@2oZ,[�@�� ��W�+0g5��������pg�=�"���Le����)��G@~�OP�ˣ<eV���}z���k4�ff�+#�h�G=�,�^5I����s ���2-Q�~�4)���	N�RW>�1��¡������)��Y Ӵ��\Yxn���iB�%4�4D�� �Lh��z�ld��˘(���O����#h-/"U>��tAʄ6�e���\q+�4#����Â|�߄���A��>�� �������	�A����E]�5��CL�
弬�Nozz&I7���� B�zu8�f��L�ߍA�o��8��c�px�oj�,�U�-�S�@�Ī�)慵9W=���;�-A�g�H����Nt�hBS�gm��F�Ў�x�b�W�3cƘb��I����)4�H�wg�����i]n��8�b86DDRr�Hx�6R7qx�N�h�������[)!�+99z/�n=�'�B�tz�?g�^`��ߏ��YF�i���J�<�
2p\1l�"B����l�ASt���s�r��� E�����2(������*M��]�����j���e�C�vhm��~��e�l{�N�;.,����>����WP���る��e�evi),P�]���u,AN���(#����)��j-&7�tf�7s&�Q\��G�Z?$SD�l��7X�a���#_�� 4�ƫ�hBS�������6ϷX�8T��?��_j�Fq��s��wU�@���ۭ2���K!G��e=�n����B6�#��	T6����;8sΚ����	�q	rY[$y#�a!���*u�m�ڶ�a�N`C�)X0���覃L�1�]� ���e�,I��g��ɚ�X���}�伶&�F��k{�9��׏Z���A<��&�Sѵ�Ӱ�x8�%�'�Ҙ�JDz*�Q:�Í���N.�S�d���Zk�.Q9�Ϸ�`%�6_'��[L����
H�U5�Qഭ�"�;Kࠁ�h���5Rv���aNd���%��L$@c1��r�\�#�'1˟�n_iT��Ӥ�5�!�8|[��!XD�o�y���Կ%��&�!,:�ܭ���B&�9BY�����>�Db��jy�PՌ���$�����<EAK�&�i+��ƅn�GGDhv)�g�y'n�rcU!
�(H��d7�ZA�)E�(s�dz��ش���#�����GP��G�=b�c�VD�۲ץ)��9u��o�f��f*��P��Ց��2'�8'�� -k ���~�R����Q� ���{�i���~Ou��O�g��|vN�=!���[����-��E%7�PmO[ZT��'|Vb���k%�<)�}��-��_c�Q|
"�m=�υ0!$f� �b:�BCJO�<l\����b�7����Sq�U����7i���} .�C#�z� �'�$G�������͙S���6��N. ���w��L�}��#`F�]�zj>������s�k�Q��g��Q���v=1)�{��wj���[q�D����%�S��̮܊�(3�k����M�ԓ���퍍sCT}�.v���[����f��4kr�Ljy�OI�O�D��:-�"�$'���e�)�%��q8��7.>��*	AZf`[��7��������L��'g�3����׉y�"�,�ީL8%y���uK��n���߶q�e��e�Q_��0�U0eD|6��[-�0i	��i���^�ʱNC7��#@�}ˊM�2�/N*�b4,!";*Y_Q�|�A�$��E"!.?�)���ӵ����fv�RJ�&P�����-˓T��]��#ȣ*������Lo�q�0-j"��46�?�Uw:bMs�������3�']=v,u�Ķ�7�|�Gz�!�M����U�,�0�h�ةV���E��NIJ޳�h(���ޒ��3�d�A���]���3���6噾�����H��u��ҍL=��D0D�٢�ӯ�Ӭ�v����-������@��G���'gO�8 涽�v���H}بa0n�{4�����-��$ax<����oA���.�^n�Wa/�� /@�<�a�ށV���[|;l��t%"a����YY. *"mƎl�d��`�cl�j.����5�ʤJ<�|�����ƹ�7��}��z Č�������{�-�и�t�&6Y���i[Q�T���%s���i��J����"L��WL��a�\��A���r�'�x�}�-�8�N���C��q�D]ie;n��2��4��k`�����հ�a*B9�-�2S�!P��O�K�8XӬ��h>�D����]�EfM����F�~^<D�VV%Fj�i*2ڀ���E��x)٠Ld�������|�
�u'U8����W�=<�R"��<��q�1ut*�Q��?Dc[�$�ZJ���.Qr������T�������W/f������biw�?0�GD#f�i��%�"E �u�В4��0�U!�._ ��|>�b����RR�lWk�-�Z��Kva��>FcdT����*C��Ik�?55>>�����"ƞn@��4i7.Eʄoq�qn��4L�2|�n�]#,S�"��[�˯bK�S�Q���\n���@�<� ��Wp�`�EJ���^��l��������zƏG�zֲ�6Q�^�+*���2�/��|�')��?�Y�ʧx�u�N����0�#)!8M �ħ�bM�&����8�z$�z�d7����=;���`EaQ����TԠAkO()[)����n˃O��5ꡠ��Ed]�k���
��m�9��ʆ�Q�����YqPNd�t����|~��{Q�k�ѹ�ǎH�bɳ�ȥ��)Tw�(tQ����S5���|N������땺g�lh�.G�~��-���{s������^�aD���V=F�9<�����No�kJ��x3#�`�^ahQZ��(�!d�X�v�d���9�h�`<����Z�Y#"Eqw-����W>bdR6a3�\�-E;�N0�}ʼCe��S�Ug�z�8��c���k�] �kZ<��L���U� � #;��IUQ���2��*�0������4��o~�&�e��6�����_��i�ڐ�u1��÷��� k�Ѓ��(@�N�X)�I��+m���Z�ջg�������%�P6�`i��r�V�F^�hm��_�aE�o�MCJ�vk"�l\�L�6��79�[�Sئa6?�[�[J�U�݌�Ƿ5���
�Ik��f������;++����#�"��q`���s���N���&�b����ʢ�k!�T��C�?ocq�Y��Փ�T��1(�>��'�v��]���\
$��X_�Q����̕������iO�2%0����4O�01��?~�h��s��H���re�"�9ݩ��/ܓ�&���e�u-����c�dA���uQ��������@��@�6�QZc(k7P{���/��,�yv�Y�ҹ�4
���oI�_�[� 4��f�%������?������O-�W��>"}2f6m �����F4U�p���c��SlO�;q�[g#�ֳ��,��'D�3 �Ⱦ�tM͇u̻Ge��Br�Y��Xɶ�T���v/�O��:�6Ol�2�LKhq4z�����w�2��w�7oZpފ����,�P�M��>���TK���
��D[VJC�C��<s~�%qi������AV�d��;[η%x��x������n�ڱ�8�3�`��ۄu���Q�_'�$�R���|����~�o��Bԙ۫��M5 �-b���L+�Pwi�"�������#�@�J9��n�N��[ƒ{�w���i<o*۬>�1Ѝb	G# �c��'ȢJwUc3��B��=�b�=q�R�Y}�������ǘ���]����l��N�}���La_eGi�bszL�Ԣo����=sB���,�kcR���O������l�L#�C�bu���׈��uv���2�##���z�]u�p#�wg+{�d.P�&i����x�[���h�m����"uJ�5��R�k"�<�Cw�����u{�F���ʪ�t>w�L��y�4�(�i�p�%S z�,.�qOB�ѓ�PH/5�85��L3��I|��A��v�L#��M���M��N6
�+�=��G,6ʀ͞C��ay�s��0,ݖ�AdB�(�d��U)��k/}���a��SC���/�g���:�%����&�M�v0��M~3Bd颪�	o����H����ζ�����s�LS�(GkŉK�$�@���ߘ�5c'��rqԞG�4PFS���K���&O9�/5%�g��I�I<L�FE��>��C�:�Y���_��6�-��B�B�E��dE)����/�� �G;M���T��Z���d�P5�1�Uj ��k�2Yž�e��D� �k'�O�S{���w�|CF��Rj��R�����͠:s�!�r�;�Pk>,��om=T���7��LH��$�[n�0 ��h�����݇�y�/dKi  ���v|�v���/Az `��k�b��gG:q����A�U9H&�p3��%H8�Rst��3�Cc�O"{4���/�*vZg��-ϳ���?���.�����|
yց~�<�|��=�'Q7���N�L/��-�
R�d%sl`Q�
��}�^ԂLHs+�a���ݖ�si1�>�t��;�N=�kᣬZ��F������7�G��Jm1(��ӽ&���<�/`�ܒ��sE(ɾ�8�+�ݨ��	�U�ɧj��0̯[l�۴M��G,Vq�?�L�/�iR��hk�����"�fe�����tr3K�vm	YYG��
x�O��C<^�9�.8�Yv�&� v�����
!g� R1NId�� ˪u���'#>�}c[�+{١>Jm��]&����Wi���8��w֙��˟%H��`<s+��#A��ћ.�飁K{�!ʤQ��Z@ت-�N$��O%j��K���:���}ei��Q+p�t�2ƞ�)��p��+&N*�#�"	Ѹ�Yo�74�^P�8S&,Q'��GĂY�����>(qݵw?P�L�P�x�H�EXlxVHYEB    fa00    16c0f����� 4yh�lz����(lV�4�|��� ��3`����j��� 
O�5"$�an ����Ѕ��M{_�,�����?Ѵ	�q
����l!�[9�9��:l6�i���ճ�E�<^y��k�$Wx���^~�-�s?蜿.�}Ea&a��P�@������K�;]Ot\r���(`�r�h�3�Z��V�7�O��uT����)����}��] �v��}ΫG1�XCK4�ً�8�]�c�֕H�8�|��>�B�&X�������'(����UֻG�B�Rm�$*[h�a�l$R�9r�`{��bL2�����3H���*�8�M�fkbc9w^ܣ���9�.b����X�xw���Bb7&��崙E�#��^f���޹��ޒ�qN�����-�.q��4���^1\H��-
�t54��j��1[��#C��̻���aE���4{��)21��l�I�4�.��M�ix�DH�T*��L� q�ư+�nq@�+O����0�k�������`p�_.��\��RYl{��R�V�}��6��b^F#���#e���f�J	�� Q��y|�{>���?x�g���ūOM�)z��7dt|(������(�{�������s���%���w���6S�0����a� �̅k��]��'܁���F��Rʛ�b�J�lX���IW�����H�.�?I�q��|Yg�E��rѪ��Q)tk�& .!��:��؎����.�/ueeġr�<�����$N_�>��{������#����#�U�O�[H+��}u����-���,i����D� Y&+׆Lp�ga.)�RI�x�.�çˢ�5t\��H���f'�:��M&�����rJr���B _��7��vP�3΋.lB졇?�C�@&vʹ*����D�dS�c�"Q�%§�!8����X7�,��y�&kL�}F����f�v�F�g���&nSP"�MbY����g�}�v���xVbN����4Q���;T n���
����Q4���6��K��@Eь�}��ݤ�L�w&����>*oV�y��������ղ��C7�BN3�X|�|u!�i����-g7Y�s6�EN't��f�<���}c���\��>�$|��5#<�]���n�$�}�`�&q�����n�������uS
�b����ʬ��v^{��(�z�f��&����Y�SQ�I�����8�ѥ:��;������Y�/s�Hk˄�>�f�G��?�p+��84PN�G�@�����K��<r�(�vQ/b���@��]��+r����Z����0��Y�55pIO8w�����f �#)0�ZL6�3>qWe�LA�%��[ja�#�j�A}�f�XjM��Jv0�-#��w�=�ŵL����F�)?��psU3�r0E�;zCu�U�]�X/�X����m����~GY��j��qg����F+=�f��GK�pD�v�C�<L�73�*�A��!��e2�
�~:`��.07Ɉ��)��]]�6{��̪����=и�,�L�r�ܱ�u$��J�Ӏ��s���ʦ����6
��Ϯ�S[֩|E+ n�}���*�	g�t�}�6���B#��N۬�@]z���x��̲�]� a���V&�_t[��Y(�D���+$_�J�h�XqJ�'��eg�kc鐵��!�^r���7߂��7��k�V�aqᇫ� ���M���~r�����1��v��m�Lp^}�(T�����V
Q�KF����-�}����S����е��XX���)V�<x�!2�ڭ�.R \7��8��zYM�"#��'�J���3=�������Dɠg�3��.�\,�!>�l�jM|�-�ә=P?��$`�Yi���Ӛ&��>\�5���ИƋ�%ъo&'\E��v��4�
N�]��fMIJ����79����-�fRWM�^�4A<���n��ЍO#W�!��j?b	<��CRT�F!T���陗?��6_�㏐чt�m�Ht'o6�W�W>�\�T�=�7�I�~��st$l��R��"�v�P�(m��Zx��L⨎b����o��G�����a��7��������;��-륯μ�8Kj��Ը��]��<W���cp�1����߫�!vGvźU����n�	�oٖ�k,ec$��"�D�.�a�9u��PFLӕ2<@ve�p�2BP�����W$��=OH�C�#Q�)&I����d� ��I����,�5�ˌ���,#L�b��jB.`��t;r�i�x�����d�@����ř��3.���Sat�_���{��1a�F"�`�wJ��$���$�9F�	R�[6/��n�R-u/�^G�U��r/�@���G���P�c��N�7_{S#5}9��JU��X�0g�;X刳�������.��7��#����>��O^�I�i��b���Oշ���s	��ǥ��!�LX ��(�$O�1/�(�E�����bȕ�o�����ZgV�;nI_{�p�R��#W:�ˣ����HJ�֦,{R���i����kf�H_�R���NH�-�' �d}�!��]���.�2=�ӧYW�����F�P�ʄ��pTIѝ~$IY[$̖�S����g-�Eh�˶��I���w�%}��:����{*������8�mU!�^r���[	Q��e���L�F�wf�ÂL�;�����YE����/4�:D���J�P Z���4�J������"�-@ݎL����`��ɫ�i*�sII
����4<�>fW!Q��&�!��S{�Y��@z'em�@�TA�%����#�t��+���ۉ��*�u�^�@� �sb�BAG�����;��o,'��,����Ym(�͔&Ӹ��:a��JV%#�#���l:�7^�tMR��}����A����}��E4T/k0HC�KUS̺���H���NBe��;�����yW�Laq:�X�HB,�~t<IO�5��P���C7� nz���*�k5��X�Ɨ�6s8���x:��\i��n0$�L���C�K��5~H3���'�2�"v�.�/6�*K���=��_h���E�>�tj��R�ssǣ��~f�|��C(-$Kv*��-�wr|��[�6h�H_�h���:�ӄ�#��xɇ��~��􄨨�ݽV*^��d���^�?�t?H?(�BU��Xd���r8�w�zn�t�V�t�= PLPj���Y{�"ˉ�Ȑ��K�O3��IQuޘ�Y�ƴ�D3ڕ8V�WM#���'j�r�ه��,�?�P��ts|.?*����:�S�� [��cZe�s�6Lg*�A@�3]�����0�i����
�PU�[�?�39�B�[�O�����z�sJ�
[xcy	���4���C���9�m\ge�	��ic"���4����
�����d��H�ߌZs�v6l����솙��ea���跖}H����P�K�MW��ޘ�>�w��դcJ���� D�w�B��t'����t�ƅ��(�s
��* �Uc�I�3 �&'��d�&��ơ��˹�s����m(��O�@}����0/�7(��>m�ޒ�l�)5�;� �9������<;�y��;�9^��#���w�B��M(�rrk�b�[���WҚu���X��eƞ�H�$UOw$��ÔU	/�.&O��@��h;Db�D~���0�%��Ѷ��S9�h���uj�%�vJ�Xkѭt�`6�، }q2N���x�;��P����&9�jf�)������Ě��S�xη�c�P��ܚ_�V�����Y�E��%��[�,��2���@>A��v_E�v-��G��ź*:G�+mi�#Q��ϟv�Nt4]��(�.�\w�JȜ�0?ڸ��:u4���v���HĄ�Y�~�'J:��л�������S]7�'o��A�1�A�%d��H�;��N�P��׳E��[�b�CL=ǜ����5���}�E� m����z�kKs�4� �`������Z�UtR2'�������-]�q��$��� j��Ni ��χ�4� �bGc�@�9�6#�����A(�ړ���6��	���k�Ө�,��nd��E�W�Q̃1���TW˶0������]��VnVhgB
��+��ō�� M�ɻ���;����JNmk�pJ}��=[&[���H�s�0X�Z���v,��B��:h;,�l]��+[-��W�@� DxǸ��KE4*�c��<*��VC���R��q*�b��_ F�3��f%c(��\|o�v�N�gFE���{��_n�������L�IZ�N�e��d�VP��m{m����vk��+�Z��GǤ�^(	�#��}0bs5x0~�@��_:Ayz�۞e��Fc�*�H�f��ᙽ47�J��M���.)�������/eq��k|�DI���b��R�����0���\�_�F�o-Y~���������
0�+���M�m��Q�G��v�Hؤ�]�=�N|�0�A�'��[����4��/8;�5 (��{��!���@�#�W�h��K�)o+�tb�u{L���a㠳�Ѣ\)�DR�O.%�A�.%4�C�ޅ���^1���M�u�FA���1^�^޵B��t�7!�i�*���8L���v.|�����#y��*���a&�L? �Q��dn#��?^���]F�juπ+��+�`1�����CSD���6���{_���t��0�`jn7��{�t�MJ_Y���_ Qk8�P#��0�RDu/~����XLd��͆y��o�.\�E|ogzs?�4рO�T��މ�;�p�����F�L"�\	�a�1^��m�+#F0�����JP�J�(Sv��d��)~����)#�efA��f<�=�}�#;�g����/�Δ>����a��-�=5汉�'i�x@�m�t. -hc���l��*������ ��AWK�����}T�������z�[Llh��B\�n�!���j��׉e��'f_eu0���ܺ��N�o��"�]|Y,�ER_cwa��:6�{Lj�8S�N
�S�{��$\��x))�����}߀�9Z�S����oz�Q��c�m��/�8e(�&"�YZ�F-�R�t�,R*�ۅ�c��S=Ĕ�>�LS-�?m��a�
G��N�AY�1�Fq�$��ߓ�=41K����)�3]�	����T|00nA��c|?w�5��8�c���&��+����|W�j�?D�<�{�{������?w��:yf�v;з���n��/
�u����RE=�%�j�)��ٞmʯR�b��RT��s��׊9މ�M��x�ˏzo�� �΅G��G��c�������������SQ�)TϪ�hnL�p��� �N�b���x��� ԜB߉�W���r�ޚ$s�'k���ܝѥl�kps,ˮ�Ѓ���cOf�NT�PQ�L��ОN��, �E�(ہ�T�3dS�|�s_ܫ���_����X*���-�z�Ti�y5m�i|�]����BW��3����gPܑ��
���H�D�XY2!���
���?�����vT3/B���7ǎ�:xe�#^��נ�T������[���ĵ�E�I���z�v�4��/���B�	�)BuJE �<
ڈS�h��Knײk�ui#����i"�Lm��f̧s1��̌iQ�l �9Uzȫ%י�9�(	���,�2�p������Y��]DC.h��*LQe�0��߹^\XlxVHYEB    fa00    1740���5�#U@8��H�q s:g��{g�n,��P�v�~���\�H��`[�g0
2����a0���E'�%(���]��~�R"�:q�7��fqǹ�>2YF���M���w����H/7���f�i�a�a�˹�XWE$K�1¼o`�ƻ�����,�d�����\��W�?}2�� ή��������A6X��[���5�nk���s�s��_v�0�U�pG��|2�MM<ś��Y����dX��h���5��a����[?�����2Ź�e
QzČ TJ�h�i:��y�������V�췖2�'Eiy�$���e�)�����p�j��q3d��;��I�i'vB 1й�G���;uGY�B�l��KG�s����=H�r�Qf4���#�l�V���Q�|�Q�_i���R�8\�^�e��V�����gI�l1���Y��L]JT�a�xC�|�J/{��&(��e����Û��X���ܜ؏�����կ�I5�Uذ~x��p��$�47b�K����`�T��P�VA)��E\u�A$�c}��$�庴bv�LS��� [�O�}��B�bn�P�6?j5��T. ��z�l�����K@,��8����d+��_�E���G�gG<�^b�I)D/�z6&�pqJ(��ŏzvɅ�;1O��� ���-LX���ZA�0��W��0}�/�1�x$�>^`�p�[�0��Ǔ�Nֈ٭}%]<G�Z�C�Qk؂&�@���
��r��y	��#�V��4��'�A+�n�k�F���F���u��4�'��I����|j�<c����i�@e��Qh >�e�����A+"0�oE.-GٲR$���ނV@5��l��U�u�e�'��h��a���j�����Y+HD�B,���/�A��MTͻV0b���	8 ��� �%�be���3j!�#p�o�L�|�Q��8s�ҫČ}^��1
��ǯ��8'���n�� eхhx��y���D�ʕ6�E�O��_i.�S=E)��ԍ2�	��B˽>��˾bܸ�E(J/iT��7$�ٖA�7���{�~�}��^Y$��^I��+��)rj��u��y�$�	|34������~��<e<���t�`Gȴ�h���A�8��H� x Aq�_=/JB��/�B�'�J�x����GEV���4TZ	���+F �����'xFT����
ǘ!#ʿ�T��xgH�Ip�>[I� �xrrN����MU��4�P�8"3�Y��q��]k��So�	�qI4�8�01�w~��P���ɥ4sC�����r�=�Qg�	3�Ȑ���x옉��jS���.�r��骇�R��Û�jƩ�-���F��&W|I��ۙ�wN�ޥ��G짐���v 98x)Q}]�%�5�X�˦��nv����@�޲ea��
�o\J��R��"b?*�r���#�~+Z��P|�ȍ^�bC���o���+�4�� �ѾZ�v��}#3�t	�X8nLeb��v8x����L�������헫�˩������Yl����_��W�o��G�4�Ŋ��w�%h�����lGco� �˖�J�gu��*���ޖB�UHB����R���U	@��{�nr��29�'U��M�'�ܚ�-��vM�$�~�yZ���z&ǣ�G��@��|f��ʄ5��a�͙C��TY4e�F����>N!%r��A�0�Erp!�D�Ԭ�P#�����@��N-����������"C7�6���� "HL������<�{��q�w?�=�C1�Î��v��a��R�6wCx�Yt�7X�~��HTb��$zޘ{�=���:D4R��]�YUY��AT���̤��|����h�J��3�/\/FB�����hW=(���WrD��X�R���n������V6��-#-6-X��٦�['����ߗP��t9t]fif_@�c}0��zF��DY�x���$Mܤ�Ϳ���?��s���t�\r�Eu�"IX4T\e`�6�p�\���5<�p.�t�`�ٴ��A�q���~�mo�[��B�F�%^r���g�����}�⬆�Џe�h;lNau��-��
���ĐA�F]�堻�zѺKB�y�i�g�`�&�г[z�K)����ǹ ���J���k �(4#a��NV�l�4�=#�#f��Gve3>xc`���/���\���_Q�l�H�o�u/���@_)�c)�ǿ������^���X���
gj�g$����-��.[��q�k�]�j�ɂ�r�x�t�,�B��){���NF���QJ5o��V���X��l���Z��Ι[	n`�[��N��zX��t4M�xY�$�տ��Wb)fOi���b�ս����$��W�����ld���(�0�w_P5�Ċ��Q�6>�:)�������tV]z��O�ޛm;�ܕRZ�8{S�����r�܁3I�0��[i:�&����fYX#�s��>4�$D[�.��܉��k
sA��S+��,��~Z�u���������D3�5�����{^�<�����܍�D&��1��b���ݓ3O�=�Q��Z�}'�\Wf>��ɝG���jn�_'�	C�m,[�qW=K/`�t��s�?{���J1M�����ҋ��h>yL9g��+P|� ���� ���M�$&r���p��h-Օ�W��/�3�v��oZ���k�e$7�3'����%ؔ����-L�|O��?	쯥�+?��O���Zj��f�����Q�6�X��X�[�[���~P4��5��l�<�$z� �&G�@r�1�v-�HC�6
�[JbE0�g�Vhh��#d��u����ۺ-�_H(܉[�����F����1.*0.94�a5�k|Z��>�ή@�zC&'!sF~gxi٭�ſ�vr�Ũ2�b�­�\DF2T�p�M����ȷ�]�#�� `��
)Pb_�[zэ|�OS:Ȅ�.�Z�;8�Ak��l�����D�X~V�o��C�}j�Z��ծc���S!���O*�_���.�L(���i���=�731�d�ȫ'&�����Zl��������"�ɉ�I�X+g������=� /N��	��#"f=���8OP��oQ֐�\��Ȟ%�<����iӷ}C�o�.k�WK��A�PA?���wF-K*h����a:�\.�+�v�镌=�՜�=�4������7�X2���Ա_q�~Y�iBѳ%�����ۇ�$0N�vg,�,�o�H�@,&��`����q��!��aRh�ն~�!N�M/�fznN-Y.g��qī�Uf��X?6�hj���B���kx�	�sR�U��������
v_Cd�+ct=y�ʘ<�s��7��,y�/5w`�Qg�G+���Be�}��<��䱳c&b����M/�ӟ�V�a��l���HGR�Xb\�/�5ÿ�'O�n����E����;Wߤ"lW�^���
2i���Nak�߳�^n�i��V��?S�\?������t��d	�3�f#�3[��$k��v�3Í����{_�׃���/BI��0��֣r豃����!Y�a���[M�o�<=��z?�#��+�+���	���~sv�)F8��/Tx�&��hYJ��0Di .p,��@G.�RЇlN��.��ĸ$�3/� vR�FL��F��8B��%݈۠6�p��F"��l���P`���A�%���{�ĉ�c��	�n�f���c������'.��*�(��Gaך��1��)}	cl�wK^x���O�SSr~��������K�,�����{��I�@!�9t)9_�qKC����S�shF9�:��S!��1�q�I*�m~k�x@;�yp%P8i`�3?~�η��FB���#G�TO�ip"e�Q�y�n��Z���	���K�
@4�d�N�z
.1���K.85��c�LOw�����l�g�07��ju�M�6�*ÝՖq���e�C�3�����ˇcyw��� w��W;'\������<5��}����;M2Rȍ����5�z=��Q�=L�&�!�
�#T��������֓��;	�G~Lm��=�z�nD~&BR��������&��\�e���U	꺩�jT<����2,�5kzj��R���neP3�p[4�P�;A�����'y���8WB-tv�d&��]��(T��=�:�cd�A�ȕfK�z�O��B�t��/`-")���&�w�S��-���&�_����`_=ܱ=^_5R FZG��w#9��]�k�XO�W���@����dt���"��f'$��?&�y*�t�
��>����#��_��:v*�S��P�6�B#���۠y��-H��,�Xˉ��ׁ<���#�Ƨe!O��9f+�҅Bd�[C�v�BO�ߵH���D[��av�9��Y�YJI#(=�Ax1��l*��"�@;�r��k��\c�	g Ϙga":���[�m���8g�8O]R8qEE���9���!NM����j�˩�6w� a/��EsTG �%G��V��9�e�����+���]��3ʯ<��T*���U�w899k#��`��ﱂ9�Aуh�����uR���!T������R2O�u�}!�Ac)��:�*1��\��F����?%�
�԰��;�}7i�������h��8E���	.֔c{��X�=3��N�F�x�g��/��P;v]��x��*�6���-L@(��!�G��7P���jɥ�˛a�4�ͺ^+���^ Ӿ���#M��zK�˛f�!KF��R��&�[������01�iכw�۶dԬMjl�-82�1KJ�֦��D'��5|	�%�B���	�����џ����ф�J�v�.b�[�����RCF�c?�wİ��F��s�vTm+�W�⻓1���U�Y��7.YZฮL��-B0Ԁ\Sf��q6],t�\�t{J5�ۡI�@�k��4������7�E��}<�̗��O�b��'�R�rX`�p1䚸t*La�4�eGr"�҉̑�|?pó����}���iLG�%~�/��)m=eE�uض����T��)T��KŴO�K�.�RJN��/7����R�U"��ѧ�U����7A�������& p%ot�[�����b�{���i9[_�!0��4��Dm�`�;�F@�����+E�`8�-�7�zb	��_�ǵ�#��?��3m�ڃd��T��9�Nۀ�zE�f���~�7aux�4�ea��Q��d�^n��'KK�J�����0�r�N
Fk>W����������C����U+�4�pn��	�Z¿���}�l�|�ߩ��6�Rsrϛ&�˚N	�w�c���w�#hs�?q!�+WώXFw���k���w^,4 �[\uX.༸l�qG�:C���i=Hp�PBU�N�[S�p�%c���z����Td��Z'}�͋0����;�/�;��>�O����y�J
���F/��)�h��}l��4z���9~:4�(���X�t@����h�;E;|�F����7O�_�C*�������5�1�9���h����97��Z��n�[`g�3��q�����.�֦��@�3x����x`k��3Q-�R�ّ��m�t�*$`�KnoJ�'9�٢��c�7'��3D3,���{���'��O̿��B	8��2�N+W����9�9,�F)�M  �����_�ui5^���Ѽg�	��\�ϔ�<�~���rb��}��`D1�Z.��Z���|X�e�U#�D�~JA�e���|%���d��#�����?Hxt�Ң7�[X:�m��)�9ڧ�g�p�x-��~XlxVHYEB    bf14     c60g8.���j:,�zf�`՜�l�*�1�G�@���eM6���Crj��_-�{�|�(j����j�jǖh�2��j�/-?J:y�g.'I�F�.�h;����Ig�w��W��)+Ь2���4]��v�/����n��/�W���yb$���?#,Z��eDr��#[����00O�(�]�7�h�l�����J��<ʛ���3�sW[d,t$�Q˴�zE]�A�#?9�N:Fܩdx$��8@Ѡj�%��#��n�ّ���F��������VD\���F:zj�qĪ��
w��;oZ��q�&�{;tU����9�}��q�Wi8��u�`��-gm�Q���S[�u�zc=�͔K�7l)��f������<�d|������hj�����p���usF���_�$��x.�/����C��?�7�J�ٰ���9 ���P�5�H��t�0J_��t��C@�כh�q�$��CP�
пv���H�F���)Q6�gE�	K<�+c*�&~��x0��gS�,�m��8���:�l*vy�U���|c�����"����\N(�*GU�a�`��s�W���5������q����ݦ���xQ�18�q=�?у�'k�����\����!��|���Δ��M�d����2oV~L�-��4(t�^Sx�@U�6�-ৱ2v8K�n��c�a�]��y$�av�'d�׆k�V�q�:��O���
K/M�b{����5A-G���*��v�X�@J\��P}o��<������r��yj�	�&x��sU��[�75�SW b�OaVză�3;�i=|�oE\�MJ�_
%����!�t�wF;����hHN���o��m�3Di_�J�&��m������5E��U/j���<܁��OP�w��\5�=1\�n���Vn���ֈ&�՗�]*7�~�6�M����������Z��b�G�t�3V>�zz2߅�'m!h�cɰ{�"�����i��"���N����S��'�T����ҙF6�#����>�-�W�w�v��P�f�j�ޥ1R�����m=}/��
��Lvez��|$Ϭ��;��
�V?����1?ZV�'�KkX �� S�֮��%墴�ܒn�5W!X���{dg����o�)�5�j=I���F�j���}t׉�����Kɢ��M<C�J=5B��@��`�O��O٦^l�O���t���oCWœq�y��@U<<��q�c���1�-Rr޶� z�:�׵go`Ω�y����8<b0�6T
�d���#�v"4��Y�l���V]P5l�Y�P�a�r5�sT����xw+CRg�f�(7\��>��:��곪tY��9btȁ˲����_�3ڂ�t�x1���*�U�L��)��8���!�Ǩ�&]��FY�QN��[����v�6/X	�j���m�����)9se��x����m��v��4X<�z�p�9��< hd\`�I��������|G�o��ddc#�[枧�\pT�P�ウ�%� �D5؉�u����|���e�����	��/��!������]� $�����M����}[��s�[;��|:I�C�� �"���û�(��61ɺ�c`]5�f�	\g����QƊ[L��e(��LU�F�CX[�	W�^$׋1��@�B��&6i�X;E��"��	� ���8Wmz��/OU���3F����7PN��&�J�~Ɉ^R�c��7�� Q(��h�z]�ɯE����wO�T�������� �e�^��M�}��$PV����(^�� 㜡r�UD��b;�ߤ������Fm'ҫ	����[�Y[m��l[�s�tꎡ�ǆ����'t������~`��U��׭�B�V���`bĹ����%P�&�t$ו��-#�=���O���-�"�g~�Ĳ\���F�m��NyΨt��xf�AF}𓕧eL��W�<1�/�y�� ���u�vAI�:O>�<�x5����G"$ť������Ӧ����)�K'���� ŷ�~�#����;�?y՚	�e�5�y�}?������	�fIҧ|Ak�.�_\��L��Do�';������[Y7J�t<����A��=~&x�In���#G��~�,�L��Tuڰ���=�	��}MA�)LG�@��bh�J�V�E\&j�x7&�"$GK5�[�L�@����K�S|x�.i1�q۹8}*�mI	���JOכ��n�*���n	L-j�aȱ�x���P���ʯW�	e�;��T]�	 �4����5c%��B8�6e �Q�lN�y�K'��J%����S���6�h�`i�L�9�#�Y��Juz���c�ʂ�u�
K�&�lwb[&Bv�!Q�� �-.�vD�$��d��n� 	�$�6ɳ���Kl�S:���ɓ	Y����O�bx����.�d礮���N����%_�ot�x��⟰\y�,o
åH�8���?=�V�(PE�~����kR��P�G?@��	�B����U�?�צ~O3�9������H�Cb|� �^���뽥�*��@ԟ���W�v|�����O%-��B&#�Rȭ�3��z�%��c�:A��� �1�k% _l�n�{�_�,p�d`�؋SV�r;��5�0 slcP��#��M��Ҋm���Τ����:� ���e�F�s�0�FB���@ӿR'��dʊȪ�V����l"���H�8��rJ�a���L^������S,Q/�����hCjƂ�RIo���?�%�����	�&{���h\��*�WU�KZm�,a
)���,f5���d�����z8b;}���2I�S���������l�U�dK�2�N���5��WBl��1 `��j���=���+��
������s@�p�X a�8�k���o��-f����0Ѥs��,@��Z���l�d�t:Վ�<��K��ᴠ�,M�`�����ߗn�B��jU�I����V�V_եΎ[\�H?�l��<f��p�A����hG6�៎�k Q���).�zU	=�q%� �����#x�{��	�I������Rȇi6�;��@