XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���E�➪��"͙.��KR��'�l��)�4���[�����Bi{���M�i.��������c��w��6��{Q�#ݮ$�1��B�dgS�ȟ[�Cʵ�ՠ�	n2Xn���ie~މn��.�I����BT&��9
;7- Ni��T��CdҮ�\f�����iTS�3@ �G@�C�M�ʲR�lHyϢ��?��[~�aC%C��{�^�p��9��Rp^\MŨ�8��;�G`[��g?ɯz�j�
��7��9��ؽ���j_Mk|$��kԆ�+E\ʳ�V���;,��"d�-�I &���]|y��͜�>��k�R�	%SXN�ٳx� 
�W�1�I���]�@��Tf����0��ao����y j�	��� -��F������{Y�e����(60t�]���ꇸ5�>������O�=���g~	|�w���`�ڙ���x���"�'�כ2�;-��|�oa_�y},�e4�@sH^��N���o��6K,@�9����*a����d0���n��b�9�*oG�q_/�G6���\��0���<�2�����C�X �A��M�S��U���X�:5	$4���p��'	��]���[^M@I�o�؇ѐ�׽&CKb�2K+BC����q�����# q+Άe�F9�8z�QEw���uf_�I&H�0��1�V��J��6=�!)2�Ѕ�HD��^î��x��dG����K��]�w�t������JP}�Eq��mG#���U�XlxVHYEB    fa00    1790�DO3��tW��TG�E��dI�[2�ʙ��3��X��V�a̴�V�����X��"Bd�b=b�<�����ϭ�}[�κ���@AZ��M�ٺ#��>V��K�绳�q7�5�>��]sx�4'0�;q���fD�OX�)]4hy`@y�Y��/�tj����G1f��v��ES<��y�A��Rz��m�X��_���~�o�^�
��ER�^T�P�x�cXb��h�ost��3JMP��bAf�,�:���!�̊�������RPd\�QZt$Uћ�T��Zgĉ�f��s��]3��F_p�G_gd�Tӯ�`#�>tO`*��cb5d�鮇��,����%u��r^���/�S�Ҷ>�?�V$�������QG��V彉�|q�����
�V\%}	�ը��
��e����;��7��[x���hGq�#�/Q�[���;���n,ڷ���"N��υh�� s�������	5��C���1��V��{K�J�2�J��T�_e�����J�*@)���^B��nN;��sl�9^� ܕK�k��G0��c�)}MZ��!�D��%�@���('N��c����B�~���%jUá�/�ɶ���81�T����O�t^�Ոv��%׍,,����7�(U�]�܆�v{vj����[c�R����)�~+{���Cih#�M,H�a!�(�=������,�L^<��rL�]�E+8j0M���vlD-��A⋲�QWA f�-)�^��W@�O���^�b�-���⪻;��qu�vp�G �w��1�اq3w�%��@G����Ў���G��g|��lZ׮X�NFy'Ĩ��ش%K�6�1��(F���Z��W��y��^�i�~���Z��T���.x����;���y�/�5.����9��v�/��ds����Pr'z��9&d͇T�F�������I����i8V�V(j}u,�E"}6򟋋�Op�v[�n6�)
xv���=�]Zc��5�d�i
q�\U	���kM��V����c�� ,r�N��=�x'��f�ق>C�OKB�%v��Um�iXo��v���U�l�W0H��7vv�m�TL�� ��Ig�r<;��j�������Y!���e�G��g�M[i�X�=ٖCNCGC�`2������@�0��7v�;��i!G������OK
��nӾPp%��&��$���'�+Mo��~����`Vխ-mN5�v敢M�#XW��b�{����z���hL�UGF�Y��	��Z�T~�d��� �g���Sc�/WG0!�w�k���F�i=�H�W$��rM�_=X�P��+�k�����X�>nY�:zVS�|α�4(��V��@,J�ҚT9?�(��<�B#1��B�Z��.� �C�� ��|>��u~%K�R�5�Y'n���4gg��XK�>]կ,C�l�C�6; ��:<n3���0 ƯM:s㊙#���.�Cg�k�j��@�e��N9
��rU�;���X�d*^��)���p�Ң]\��;��t%ռ۶�W��N9�P��%r��\f�"el��#�	�r�	m|��D�k0@/X5��N`}��ؿ����V�����bN����X t��CJ����jNmI7�Io&�yf9ë�_Iͳ��K=�Ǥ:�5�w-�Hh�/���~cAX_��o$N�g0��jmUZC����*�0�ض�������������~t�%���O�%���΢�u!Lc�t�Z�n���4���<�����!���.��+�G4��g�� �ɑ���Fq­viE����4��{���Ɋ/�04�@�UQxH|kXp�K���5B���"��5M�Ƈk-|��$Nⳗ����� A2�{��x/͟�vE�=�l4J�V=�}��p3���R17��k &����+;>��5���=�;�~K�����	�~d�N9��+�XC�k���46���L�q�#��[��.�Σþ���uB���U�L�Muv�� �9�N+���v[<� �aN�ט˲˴��"D)�,�4��>�a	�'��ӭ�v�y�Ƨz�3��V����S�t��S0u��]2�Ҽ�ཙ�0�����9�B|H��x�8CQ^&c��
�^U��s}1�Y��q�G�Z�N�A+��~��s�}Ί�:�C!��	���?Y4����˹6�Lm�z����gi�/���U�1��G�/��F��z�B�T�ֶ��Jfjہ���ć=.�v�G?�B%�FA�������j��%��0`S�^Ƕ���=q:�)��y�嵵�p�m�M��˭�t�������(�z�״p|h��B!>�IGvo����}y/oN���fo����z�j�m���9�f2�Dk6ȷF�"w�Ӌ�]��UٗX�v�V&����,JtS�}i�jrXO�A�;�he�o�:Y�m����%�� l���	2�A�$��
��(���Ep���Y�	��/�n*��F�8wqC}g��A�2&{szr��z6a����~=�^0��ڥ��Bt���6�a|�p�z�bv�Ik��Ԍ�B[�x�5�ŷ��+�O�e0[�f��
�' �%��0�j]U�-��S67�@�w�
�k�#���q��_I��+M� ���������-h_qQ�m����꿧�z��%����i�f��A�`�.B�����Ośw��s;I��_�e�Y����nG�d�ݍ\�='/���ߔ����5�S��A}y1�����x;o���R��p	�%����ٖ%�e��$�'�#I|�i=	�{ڻ?1`p�jr����ؐ�QER�V�J���^�Q�L�xҙ�6Qa�"`�I��]�I�R�%����)͇|T��X�]��6Iڅ��q����n���t�	�1NlvS[��hP�Ni�\M���4#��ޗ�w�J��ͶB��hF����|^38���4�����p�_����M���������5��W��
`�%�6�M�|IMN.U����
i�Qm�&�M2��Rᙁ�i�Hv��ѭ�Y)}j�$\����ʋ�g7���ps�,U�>��\6F�T7o+^,�	I���Ҿ��H�3�N�~=α�tF&���]�$!4��J��;�U��Y{"U�^	�=ϙ��Z�V���>I~:�[z��~�sAbx q�?Л�/yla�_Z�J�Ӓ�_5�`(��/쫵H����hº�7k=�i�X��ЪQ?���C?R�k�*����0|+i����^��-ɍ����wi��%K��*���!��{ص�4�� ��z1!6�C���ީ5aB#܀>-ީ������,T� �U �_��T�z��]^�ű�N�O��) �t,q*q��3p�8x�ZӁ8P�O�4�`+��^�����w�C��u6�#�VYP(���6 ���~��Vf%³����=73�$o��g���\����>���e�$ Z�`;�N~ø��Q�7?�\���&�=d��OTm+3�&����p�ɼL+,!%s�¾��=eN>���},N��U��i2�������C@��C�FH���c�ce߼���~��I�˪��TrP����x�R{�H�!`@�}�-�Cel7��[���G�qQ&[k�1��\���-�n�%q��^��T��Xz�
�������F�L����`~�@O�a�cܔg�@~�aBA&����?4�G�ϋ�/�7�]J�=L���+������59m�8o�h���`��z,����>�UR�E�:���ѩ�or3�U.��j�ΞG��=������&�G�t֖w;�PN4h�n<���O��" -������(-X-��6�C�njzZO�w�?u�rV�~���-��'4+�	r��;�w���Y��@N0��������-�I@����ܱ��*5P��p����c�a�{�$o4���l��hV1��S������!��ܪ����&u����2�<Bn?ss�͓c��9���!���(`��(���~	�P"?��K���j��Y/�d
1�>��b�~6ڒ��ޑ^G��S�l�y��r�i���n�z�B�K���Y,�q�[�&��q���9��<��-MU}�6�utP�Z��3�k-Xŝ[��5m2jbK>����`�䒘�T�p��9]��L�t����	ӶhU��th���%����t��F�+A�1���دQ~�&��'��A�-���-I��}�U�jɢ���V{�kG�E�-�~� �aD�ct/8h���M6�i��5Z�&�Dwŭ�W5X'�W1��:�È%����Jɪ��íb����xf#yWF������t<m9G�G[�RN�t��+��[��o3��ݲ�I�\2�B�:qTW�@DB�R|�?�@մ�B"tq�Rd����]�ʶ����PD��^�Y����!@�y%�$3�Z�Q�����<F��y��`�\9I&U�����P������lΑW��V��#�P$d��%P@��#6��q���پ��4f����CPds��>�-���N���Z�ى���Fo�W�G�w���p�}���<����ό��l�^�)d%o��I~���O3?��$A�xwB��$v�����"CEl��$\@ߩ#��C�#�R,��T��U��`K|6�n���j"���u�
����;[l@��Cw���6<���
 �UuÚ@[[4�w� ����u�>Aҵ�#@�f�ޢiT�G{��'������d�.���}�;s���0����<Q���y������w/=��b�JW�]J��_���*��NIs{��m�6L�
���V��V��%�w�#��=C�;3C�'c&��>�/����y��
H��Z?�����%;6��m��:�u�b�{L]8�={#�R2P(�K�r�Y�]^�55@kA!����yc$�.&z���K�����?z!~���=l�.� L���ȟ�FoIӗEP� �a|��;�8�ᡫ��B{�Z�kn�.}��o������C�/	��cg�`�k����x2G���̲Փ�����2u��KH8��R��FN����s�^��69^�rp�W��H��Sk��/A<648���^F�3 ���'EH�G�j�:��'u:�A**�_�c+��P���>y���������Kf�{�(y؝�A�����(���ϗgk�Cb��Ҙ�
��#I.i�N���.�n'X3|�h���?�ɭZjI?ɻ_�ud�
{��3�,��B��� e��ܹ��[���f�O\(7��Yo���+1W�3YR���ֆ��%�b;�An+:��ۑ���8<�w�C _%~C1�7�Sܣt̰�2k��Í2U�r!��Qx�p�����$?ri�
�N�T����^��X�*��<O�)�A%�IԊ� _F�O��{8F1�w6(�"� �ة�d��y��U��Iji�������������X��#�u�ǥ&�혿����l�<u< �3L�+Vm�݇�V��F����xTFL�/c�~q[��`���t�`Ǖّ��>�^���W�l�خ�ꔸ��2�^�BX����b��'.2���ii���O��Xon��w?�3r'���Fc����2S5&�1���pj�S�Y+͗ƊQȀk ��~4���t%��%TT�YT[�Q�Ԍ�Ԝe�v����^�p����K�mbi��̾(yT��v|� �	�!���& ��n�m��m^Ͳ��~=�v_�#�#t#�`c.�8���b�C�fӧ�o 6kM.��@����c+4$?���c�˺��a�����|��(�Mq��W��.$��Ad8	�J�,�Q�K�C(���N�q��V@�=?M=��y�����)-t$tf��P0�M}��(�.G��N�c�?�R%'��:A3�a������W�ٝ~�`��	)ʘ�[�t1�8k&�t�0y�m��7�XlxVHYEB    fa00     5d0�������_��K�GU6���b����6�]���ϲ�^̺*�c�øx�7����C����n+qߋX$�ǣHx��)���jU6K`�W�bk ��Z;���`�2ϩQ���7���	�͚HG�\��Ě��E��!"7س�����p�~h�T)+7mZc(����$� @;{�j��6� �r�C�'=�&-i0�f|I�ҐQ�o�A�����.ʧ�a���@.R�/6�1�Ў�B���Nfc��y�g����F˓��(-V�m
SGݽB��u�X2BC2�����&8��8Kh��;ȷ	4ρ�w/��쐋�H��D�BΧ���8h�|�X�ky:�W�n�HZ��=�le�ӹn�Ec5��ɝ�~:�4*�SV�x���_F��`���}@��f/m*��;��S���^�)�{��{Oq��fw;����;�즃
D�z{���&�S�,� {���WfY�˖�a����Mh�p���\�6���h:� �k�%�͡!��꘡ 1�A�t�����g^&�ak�Af��_�wM�M�.�joN���7��BH���j-��?��5	XT���\�o1=�c&���ҝdv�j+�@��M�T\�y_"݋�5m�wg������e�H���[�ޥ�/C�k�(��Rr�-��n�K�1�>L}��8�MǴ)����:�gd�� �[+�
���Rm̼�@�QIvyD��\�x���bF��y{ .{펈l@O�[G�.\�����	OwS�w�6ɬ�޿���6��bU�Fѵw�MU�tj��t���O 5�I���N��k=��q�d��"a��Vl��ι��q֞٪���I�.)6f����vsǽ������Lj�!��_>��-1W'F�L�F��6�_�!�Dr�t�2F#�fn�A�.�@t�{��p��<�dz��F���v��[��G-���ｧ��+h��7�vi�{���5��qA�"�������Z�D �ā��1�aF7�u �G&�����>x8���T1+�����؆2�������S]c���엡�?v���������$Q�Q+au>��4����.�	�)oI�:#By��q� ^KG�&i0��{�>&$�P�ܚ���� ���U-�b�Mg�)	"HzD^���,�b�k�ldx��6,vK�䅹nR�t%0��S2�e/���gI(����9*��M�L�AȂ���8�� 3��}�����Ḍ�X̩(�~��)+q�Dġ�J���G/�#����C�C{� L�]q+c���9�a�T_�W��~H���ҟ-An67U��#��)�����7�v;F,����O��^5/��Ep�F.�D��AЉ
~�1�3�{��-<�2SJĜ�2���D�Y��P���C�"�ae4#pG^��;0���-�uӾ�5��0���Y �K��^������L*>��=)XlxVHYEB    fa00     640i����J�HmJ	ã(������z�P��a���h�wy�{���?��b�k�3��ѹ�ׂ҄뱲�@-��s��A^�p8�x58�j�K�怇�|K���01*�z;��R�v�����[Z�Ok�������w���٠ۻHZ�K82wUP��l��)��獪\�Jp�!��p���tEM�Y���T)�G[j@����-P��O���́ڙ��3^� hV��v�����v���+�e�ne0�Q�ʟrߧ�����y�p�:�m�ϟÀD�#��@�f`�!)o �OɭP����=��atdA��^��[:�mXjM�mڟ�HC�|U����?eV��e��m��P���/J�P�N���k���_�,����lhO��bd�rlL����3���3T���w5�͡2ϊGЌ[�
[$YW �q��4N��� ��R�η`0�D��)K� �A�ۿ����:5����y�����E��V[��zM5r��DKd/Z�����I�I�I.�Q�	ycܦ��]ݮr\(��*��$ӓ�UE�Ik;��+9��D���f��q6�T�l��p[���0��c%�u�>�
a�XR%��s��߹0�m%�R������Z��&����MAMK~�����+d���; o���g	o�,���-�\L���*fX���敄�+��"F4�����
�����|�������8�|g�O��=M�ځ)��."_%�Rh�YoR���ެ�����4[�F�I��{;�D����+bu�.�F �#���]�,1���+uc�*��)F*���G7/��W2�e���*���J�2H�b �
<�(-"�<,$���d��p�b�Ã��рԿe�R��T}ڊ���A���N<o~\�v�
�-Ċy�a���D���	V��n\[�O���f���>#��-%��	��t������/Q�_�
�xg��Gڌ}_ْ/��)��P�|A����j�nz��[7��4z v��-��/�g�.�v<��cZ���]�WS�+��ߤ�|��qY��@.�ݓ�a���4M`�9.�L�w�i=�5�GH]�=�p)��)�`�� �8	.��`H� �G��!��㑗{hqM{�4�D��3��"%5��V�Ӎ�������!/I��6J�_1�u%�,V��ʂ��f�9m׮��0�7{+�*���[�/��J-�(��j"T��Q̀�/V�l��{�@�������F;C?�)gKEmn0��j�_���6t������T���U�!���{IX%-	�oa�b����,w��q9��y����^#�����sQq�/~�ɆBm���ƽ-1�N�?���
Y��2W%�'�XPY�z%
���{��>6P9�@$:�ڇ��e�
���0����Ijd�=5������@�����o!��@�EL���(}�z�EW��"�L�#���l��p d�`V��|�.T��qE.1�R�9ۘ��|,���E��e:�� ��*�A�
�n� ���x0U��ޗERz���M؉yO�Q��@i3<&m�j��.��C�Äam�tm��XlxVHYEB    fa00     5c0�ԧ��4[zޕȣ桩�k����
�`	;o	�&�RZd�b�T3$�4�~�Q$2#,v���$��O��(��@05�-7g-l7�`%U�ЀBz�I�����o�-�E�<%����jBé,����Z�m���v~�^��If_�3�����7��.�c��V9H�y��6�}�����q�~�t�cF����!��w�;P0�;r��NS��h����t��U��@[�"��)<5�`�uLA��atbU����6��·t�-H�GX�Th�P�����SE������r~i��ƫ5����GQ%���//)D9��d��܌ ��&9�����<��s�T��_���`]4k0�
�VY�S���&�;��Fճ+A������knr�K3 �c[3>3.�Ջ��{ϣ��l���n�b?��Y���
�}�!��g۔#B�^���̟�h�P	k9�M>���ci�h"�<O;W1h�"�%0��*0�z��0zK\��>�v�/�v�G�Bk6`�3K��	}�J�l��w�p��֌�C�BC�� !��W�u��}عę�#��!�˰"�ZU�,����6�h��d�p-P/�������o2����E�G/����AX8�E�4O�굷�!��ry��K$k�x�K�B!;�v[������%C=����w�՛�#x�|�O������#l�
f��עk��k�+B��P�t���gf��K!c���U!�)��+++�擂�amX>е��L#�J�w�>��^�2� ��i߻,�b,�:n���]���ɂ;�x9�֣? �t��b&԰`�WT��g-('E��q6�|%ř�j���t�s=)��e�]����#X���	8xD�1�L	m������4�a[(��J���)��v���is��:٦������bA(DwK�KZ�W}3�j����V8�e@���.�<�\,' ���烂T��7�]�n'��>�d���]L�W�� �\+C�����U�5�K�
'����3b�o�*R"��λ��8p(j��9�HW��y�����%S���cBП��UR�z��ro��ޤV:���T߁<z5�vNRd?�-��&A���݉Ƀ��c���/ Ief��[�5pV�����×1Ιxa�2��w�As�
O�s	��Ղ��n����$z�o�مV��xk��!�1 +p��Ԓ�Jז��q���8�OӫZQ��������ͥ��ͫ���ȥ���U�1��%���Xuu�Ѽ��']h�DQF`����Z���#U�7.g���L�F�]S�ZJ��Ә|GĶ�Rr|���
��q˂~��-��4&��۟�#T�����E�[�L��y4d�q�w�e�xZ�`��;��˗*�<e:ap�������a�D{�Lv���ƒ7�Cb�'r��p
G[��da$�יԿ�V"f{XlxVHYEB    d347     a90��a����o�����gv�Iᴟ�0}e�P�i�m�?�
N`9�|1
`��
��B�h�]
�$ K+�RX�Ӌ�^]w�q?�u�ko��7���UC{$�<�$���A��9f�i�#��B}HE���ġ�nGrl���2�фՄ�Ɓ��R� �|,&�y[��z���Ǵ򋺕p���䅅32��I�=�1L ����=+�2*Q�u�G�p�xBy�ĭ�׍<Z.�^gG&��k#ӂU ��r�ܨ�m�P�|������1Y��Y�Չ��N�^a�1�G�R��6�I���`dL�t�x����zh��EjC
��'�w]BX��0�S����t&�-��	������E�h?rnPw�VA��&KS�Y,bk��͒'�
�B;驾�)���H�p�v*��L1X�'��K�B?P���,y���n1mڳЦZCe3���-O�?�&���s��-�܅У����A�d)>焔��k,&�@�L������:W�ά��aҚ���=��L >�V3��
-����[�:��6���F�h�rm������P�򺔎u�}-�E��Z�,�6z�� ���:X���D�X���ݑVM�$�%�{�����#�5>��S��R]�Fp�g:��w=q�%f��*Iv����߼u�9�\1���.�����>n�]�'ϭUe뉥Xq�|1H!��h������H�����lF�i�O�|.���V}��鎖����0��HV��v��b�4�[`O������<4�K��5��P��.,(�Ky�RE�a[R�ϋ����ӣbU���?��Қ�r	G�%��,�y�A2�/S���Hq;��j����TH�
}q��F�ã-�oq1�Ϸ�H�>���i�Bܾ�v�������%ߕ�όj����m�]t�l��Is�<�No�`��q�Bj��_��RᐟkQ��wK�҉{�M�r�1�Mt��C�{�����t�7�q�=��c� 
����t�}?u����2�x�%ePk� ��T�RQq0��-�#�L��Zޢ��9�̂$G|̍|��]\o��G��a�pːU���2p�C���XA8��m'i1%������U��],��ܫ.��ت0TL�<�X��U��rv��|�.[��O�:eFT�7�݊2��e6�}��՚��-�Wc�s@�J����Β?�$����^���ֿ��9�:r|\x�p�������ꬁW����X��SKݝ��~E'?�8M��������)~���JL�i���B
�8`.�K�8��z�7c&sk�jwc�L�8n`dv?ȄR� RKCC��ƝZc.�Vj�&��9�%v�e�w��W��Ppr#��V�'<P+�_{�Sob�ԝ��@��t���,�>հC-�"<�D�8yY+H��j�Q��5�y�_�_��AA�n�:r ���<�	�v�F�y��7�W5�CW�
�>0�{�KC�: *�u�e����'���V����$�]��r�Z ������ώ���8J��ʢ�!M���>�`�2s'm���a��i�R(�ѷ��F�����B9�@�2F8���?�y�����q,�?,{�5~낙�({d��~�"}�NU]"��<�8�MX��عQhm��4�\ϜO�w��ۚ��I{l�W�t2��2vZ��l��7��X���gw�B�<�[GvW)��hy���68�9Y�6�����`v��6wo�R3��������q%8ˬ$x<�.Іi����Qb3�������Q�Z�J����$@2�;��S ��(�(Վ�p�u�W8��k�c�l鹪�J�^���Ne]	���/�jb�Qe�������q����ந������1�}�/蕁�[�:o+2��!�w�~L埱<�X$��1��՗�N��U�!�r^��ǸZ�K��>n �7Z>�v���_\����O2�yE<�e*R��ˍntht������lc+����2U΁��$w�
�P�#m�!��'�!��U�qEsW�m`9{�9�jRK�oK�(&����ق�e�~�YQ�!�U���~8�ǭ�f�`�8X��m>��Ez'ar�d���Ur�
U]%i5=b_�y�㸊��L�*� ��3&]+��5���A�Y���n�҅��4�'���Ы�:�7d�P�<	f�cg]�R����r�Erq�Ѣx�� �Z�
h���b����	���޽7��vX/�:�C�1L%Us譈]����uV=��TfS�I`��g3��!�2c������$#�Aj���8�C�V3y#��.��L��4���@�[M�e�+F�x��\�}�te�-Ի���#x���"C0�u��ʸ3�3����1q�m7v��$ҷ4����t�z�w7�*^6N�V�����&��l�@�ۈ)�{�Byz���'��C<��{����ΙӐ��q6�W�D.���Q�5Ugڽ�I��̉ȁ&j(�P0�v��{0�����U�z�H����#PʶQ4�g��k����}���ϤAK�0=KaK�ùK���\P�]�/a�S}C2!�����/���n��v�=DFt�!t�����
 �����D�_"f���s�#�����EN�׮3��4�fTq�Y��K��ykI�f( �upA�