----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:39:19 04/30/2020 
-- Design Name: 
-- Module Name:    Interrupt - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Interrupt is
    Port ( clk : in  STD_LOGIC;
				input : in STD_LOGIC_VECTOR(3 downto 0); 
				flag : out STD_LOGIC; 
				ISR_VECT : out STD_LOGIC_VECTOR(15 downto 0)
	 );
end Interrupt;

architecture Behavioral of Interrupt is

begin


end Behavioral;

