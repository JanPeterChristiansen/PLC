XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���/?c�V3�g��q <�t⠋��v����Y�Oewi�J�Yp�c�Q��x:2Ԧ�%̳�61%�����q���<���������j:HS�h�?e��jȸ�0H3{�+1�p��sk"IgAG���H+qs&uY�DL�bʉ �;�pD�>y����tr�^D��������tuA�!��xC��.an�>�)#������}����?���6��&��0�M��n��?�u:��>�1��.��
�.�'	�1����3�p�r�)���;ږ�$�܉(?2����~�����3�*L��'�J�5�����A���ԇ����|���*�Ά���i`���L�J�����)�*����?T�(�	�c����-��S;�.Qҧ��.�-](dM�pf����݋�z�}�X��6��gg��D�ԉa�/'��SN���_#�R y���F��m1��D�١����<������C3�<�K�*�]fp�?�Q�&t�ѽ�E�{��b=W�ɘ��A>���$3��hl���8�I
�2�%��V+����U��N�d+�����-l��R� �ff�� �#u��������K�`��z��;��#��/w	 &�f+�ZD9���`N�I�ꤠ'�:��<���7$:���ې}�f\";�j5��W�?Wsˎ�r675�A{�ʴU)�<5�� %*:-�Y�� <y�Q�ܜ�,q��t8ȝ����	%�PЋ���PXlxVHYEB    fa00    2d60<%P�� �N��o}gW���������1�������HT��='�[j �[��D�M�s�z>n2`�uߘ!�ƺ�K����(>�vF��O�@�!U�B 0I�HCMA�,L��:��5H�=+���1(f���i�fv;D��"r��B5���}��`U�#��i-�̍�Th���#;J$���s= :#zN��,N@�\c��_&H��SE{ �κ��&�&-h'Op�>��\��D��1����j=z��Ұ n"�i8R]Տ���L���%��яrL�CSEp#kVa.dr���S�y�}��r��*9b��z���ftg�F�m��10u��ھM>J��p(�3@'�W���j{���62����y���d�U�G;�xP�g(�Փ��6��B�'���
�M�q ;
p���_)��tt_G����լ;�O
IMiaI|�R6�<�J�t���|$s0��e��&�RXh��(��١0#��kr�8`���<rܢR����i���㾢�[Cp��K����@4Y���WJkh��R\����A�-����o�cG�������R��;Ԇ��G�G;AY�)7[a7��s�񞵵�Z1*"�	�"ȟn����%�Jʜ}}<Yew(?p`�}j,Q��d0��&2�i�^�(�~���v�iv3�X�<!A��������[�_�i�X4[��Β.�6����R5E�ȏ�Xk?/ڟ�AK��S����A�ʦ^����uzr�v�w�jȺ����Q(%ĭ���V�"���5��H�sY�F�
[9Ab�����(*��`S�i�X�PjQ�΀�"Xm"7�?'��I0Z�T ����q�c3z���.k�2cȇԼ�����9aur�f�&Tɩ��Y��&�iZ���y�cfǔ�g)L$�n�OS�����ĕ�����5[7W���ٞ�}mT�F�T�Ǆ�=����e-��G`fAR�N�0�G RQt������)*�CYlN�cԏw�|���5[��#�����1�6?K+�T��dN�}&G�LCӞ`�,_�\��J���ɳ�U&��gfXY4&����%��A76�@�LY�����|/;�e�%�tŃ����Y�S��޹f���'fb#"�k��!�
�����ŵX0_�F��C���<˱j�#�����tD����7���8����e�?-Cw�������)�t��ޗ���-��fbp	���Ϩ�D����Sg�'�Y�k%��k(hս*�?J�o�CÁK���lJ]����Z� 5ȓw�Nt<�F��"EF�d�F��(r����.�<$�^|���|��Jv���7�r	܍��;�{�ꃞ4S���#+v$)z���4�~�Ά����g��<���%a/��ak��h�fj���Pc��sx_?K.#������Z��6\!�c��E(B��js<\����s���d}�{��Ɠ�s'L9j8-A�v�����l��JJY��k��IR�K�YN>��6?A6�h7�3�t�pI煫wV�T��w�bv���a��F�U�~Hr���<�a���6SL�x�i/�؉�g�s@1l�Ձ*���E�ͻ������DtI��ѕ�jN��G6'�b|��DW�"�}�=%�@�#hl��o��;�k�fa�YD������N�i��fF�giߖ��/� �U�xS4�1�+�z�m������~8�C恉�4s��%��"8��a�Y
��|�\��r�%V��;0�u����0�q����[.&h
i�uIN�<_[2$���������?�Qdx6�J�nʪ�:bb���Ǉ����~ĥ�!��Y�
��zR�J�8��K>1���uZ}��d�1=����(_qJ�n�.�b��*A5���PhF,�jv=:̈gna�<��y�&0j$�V�V~�T���*m�?s!�.v��RQ>'��?�7}���rQ��Ɔ>}��}���O�M�j^���Y�^�z%>������x�+�B\��b���%��v��DZ�S!��kH��%�ع�$�D��x�Wo�,\V%;@�����z ��L@d����,_��,zL0��o�yW����Z��#��R���#��k�c�n��_��ξȭ�%�H��~Cڦ��ն���,o,���	N�cB�ϽŊ�Fx���'Ri["�O��͒�9W=5z��Z��Ho���p��[�� 6�[J]�*\�u��Dd� ��O�T��D�F6~��0� sW]fX�-�5X��~�&07{Ry���X/7Q$�������Ɲ��z������ԖՐ�=���v�۫s ��Do��	#y�-;���+��n�`��gԤ7˱y�wo���;]>�.XS�_|;5&��U��~{��
Q �S�#0>��(�܉5�ꤺꨗ�&��P8�@	���q��[�a������ע-����~�cf���S]Ɠ�^Q}�-0^�ն�h����~`C���đ)@��!sX+�\BZ�*�YK��@��;#J��om׏�c�'��	�'�q�@�9%Qz��Ȼb��՝�0c�E���R�?D�8��A��qS�����ї$�Q��x�H��ߕ__��@����˫�c���ƞ0J:Y���(̿�u���y8�$��G����x�D���+ ��0-��������~���iЉQ7ʲ=e���h��J�(Ko�5@b(���O:�A�#]�s]���0,3m$�RZJz9�T�7�mL�����?����g8��E�v1:����r�'���D�ƟE�T�.k���?��㨩��m*��z�"E�����!mI3����Q����P�,k7���{|��AtJ:�|�aa��!ú)9�j��Դz���E���ғ���b�>�jч�on�-�?+�K��F��ˎW��(���ᘙ$����кף45Z�����v(���x�,0b��:�Wĭ���͎Ц��_ȿ���\����h�'�3+JzcHL��Tj��e���mP�jo�k#��/~��Q��E���|�;'mU���eI6��m(a	���D����� o�F=�J��Km]�ʽ��!�.g�滨��'WӺ�@n4�^���,-_�y�#1��NŖؗ�a�*5�ZQWl�E�+�kS����A�@�{���R ;�bG����r3��_"�7��[F~��J���H�W\���%�C7��5EX����\"t+�kR�XN}��?nn���v�J8@�`�mq��d�qMn ��Q�������t��p>h�\�Hy���ǚb��	UHڻ�~�a5��
���/����t��g�G�^p/��1�5wU�S,�m�/Lj������!Ym�C�+��9 ���%Tͪ���i�)[� �2C�������� Ð��H�ڶ~w��Z�#A)�����gS��A�!_ֈ���3�Lw�h���X���h6l��%ɝ&�V��-�m^X�:	�G����� 0���ʘ���J��ہLqpb[B���*<`��6���k�Ï��˅�SQ�ױ�8\�n}.�7`�}�UNz��͡��*��1�,�����������CpLN^5�e.�1��Z��S�}r���U�Y�(>j���F�����u�g��'����w>k.7KTj|�n��*���G~� ����ګ�z�^�va6��<*/�Tn:h�%3�z�n;EY�lL�;9�.~}�Yy)�|�Ж��L��d]�TZ|�|�H����������v5Ɠ��L;��4�~�|��ȹ�����9���B��!7-@y�3�N��ڮYby˵%f&mct�Q<�Mi�})ܣ6r���h���T�7�h�����2 ���V���S��t�>�Ƨ�3U@�:�h��$Ҕ}�� :�2v�ie?�\3P��dKq�9��hj�� Y���O���m�p���虏Jץ黎��.V�t��	R�+�[ٙ����#��<eX�w��*�/}?;�;B������	<����C� bIL�H.�A�.k�v�n���΋Ƭyc����j�;hV���M�1]�%waH��\J1�Ii��U�B� �2-/_�Zo�����,"J�=c�)��|�ki˽���kbH��a�yrX�*s�d�e�ӻ3·��8�r��BJ�#�඘Sd6IR=�WM��aewa.݉�2���o��f�E\ǮI$�hŭ�<cG�珕�5�[�O�Zxɣ�ͼ�L�W�]۝M���k�q(����8�G[�u�P������ �"��(��b�^N�,�k>	lt�*|E������e�Uj���E�Պ;\�� �����´�n���/�/�=B�Ya�&��&"���ή�yo��5���3��KU��j��3)�R��<�N�<W����4e������P䚐��˞�F�̫�/�T\P�w�`�~�@��jWޫ�FD����Tr>�9r�@ۍ�ݥ8HR�F0;]�ag���B��l��N�_-MQnq~h��'�������
�X!š��nl\8��bz-(�//����~��"���d.���Y��"�(9��c ���&�6!_�C*!���|�{5��wa���4��Ę�N�q�1��Ɗ���n�� UH:�q�&r���5?��E�Ox�� �/�rbF�`64	6��ָ
\�T4���������ć�g6¦�'����y6-�ē�46���bkl��� w�4���ɼ�l�|����`��,�2�2	�����a�ق�e ��k��!Ne���卧}d+�8H�=�(B���p<u�:���Ch9j<&��=�(���׭�t�7�Pک�~(R?/��>��Z2%�v�����6��� �y����!�e� �{a_cp�+�M����Ϩ��W��e1璘�A����w�v���@f���8���M�+��a�W�PC־��ؽ����q8�6`����a�Q�a2\��"]�,)�]@X�q�������fC:�w/�Ś_&�n@�$��5��;,+�u"����C��\$�9&����WCc&"b�_F�{<�Q��=�WѮ��B'��b�Zb�H{8�Q������|�	�ɞ�b���M�Ka�`��i�5IV��w0�j�{�k� 'ĉ��>��b8�������[#������4���
�L���Z�O�A��u2����>ޭ̬e�`���q�2$4�u&V�{�[=16��X�V�D�b��VJ�����M�ک�]i$��)�.w��K�C�AH�#�����]�qΔK>�D~����J�H�]�u���*��������dY���t�呠�������ߵn��o���޾�u2{�a+�Qu���ﶣ�ȅ�BM<��/`����1��3�I���-�Iw�u��-��hК!ϼ�u�Q��u�������.�"R�Աa��odh�ѡ먳��=K_e6Zs4�O�М)t��$"����ч����H;8U�����[ڻ�*���?��7�����+�ZݧJ0%���X����aϥ�0��*���taR�4�ĘQ��6��%S�_���.�G/PtE8Ֆ�7�i6lRB�"?���è��\L�oy�v8���Ł�_�������p(t��޿�X��<"��6��d��u�֒��eN�k&��̃mW���\��dj�Ĝߨ�+K�,7��U^T/T�]͏b��K�-�'Q�k/n��r�}B�B�b�>"��z_"[�������D�O�Z(��3��� 6�s-�ن���Q%�$q�l?݀)�܇4���-PNf�?m��}N� \��|�p�����x��X먐����;#�������v�����6 ��M���G�(�\�?=�S	tXZt���{�0>W��l��N����[N���\�$ǶJ �u8�p���uy���I�ٚ��4�(��d����������q=Ӑ���H #�o�չ�8��~�i������0G�R���w<�0�,�����,�[�30+��p��?��J�PGIN����3=��Bv%�aJ֯����˄����f���D�x��i��Gv���J�7�ß	%��,I�bS;���o��Ja��$n�_�f��(=v�SV��y�!k�X��%=�Ɛ~_����{yeܨ��h�S%�i׳�v#0��}"���l쥂�5��?�yG�Zz~�����ai�B� q��1؟�U/)�J��Ml"��̡N�ibB<ij� ����������U�,���q�8G��� -�fvvE��䘉��!�Ω�ӂ��+�a�T�o�Y��	�C�i�4�
1�1�����0Н�5yr��e7b�7����ym�sG�����f��[ָ �?���HQ$Ke��v�X�fe�!څ�z�M��&r>Ֆ���M�;6rZ*�;���c��R����"ש����5�N6hꅣA -(�2���]�*�ĠP˻.i�{�%���gh�-ɔ;�i��	�~PYm���(a�1sUd�+��"���ٻ�Z]���h�j�Nt���P8�	�L��#E	�����Z<��?+�3t�aQA_>��}
��bBt�KJ.�7]�+7y.cu�#�;�;uy���c������Չ�7H`k7̳���Ť�d����S<ν�U)M��')`�2��D�����I�d+�Gc(h�/3�
:
�������������l�<�̞E��o�g��70��)>9���E��P}@M�b���L2g��q�]e��+(���vT�r=�r`��ƥˤ�G���SA��-n?�����n?������hQ�@8�tݠX�h����j�`��w���.���$FQ�R4^
�����2����0���ő���F��@г1a��6c�0ת;b������ �4��P����+��I��~�maN?l�Eк<���XUQ���I�J�-�`H��dn�􋵀�3��H/YB���>˯1����֕�`��~���2V�Mc5��͹o������$k/}n�G(�LI+tT��݆Y�/S�	���w����Y�u������|� �+�D$��1�J�b{eI��q���p��N�VJ%2������[Eu����:�àg&)W` f��%u��vG�Lx�!�tM?m�b�}	A��ֵ�1��i/򼳒��ЉM��P�YU��H5h^�?��Sr�#�(cK~I�ע2QP��'�)�ÑA>����Z/vv�p^��پl�wid��L�q�5$��
���A��0�̺��YJCj�`���g�>��0;=I���L|���Ԩʵ7�rk�')��^��k�W�!���>��Md���>�p7u��>�B�K0'[�����l���0�u����q�}}U�$y۰�������A�BQ�~�4d��|�ɵ!��Ԕ#�>��)ڜ��9\��0�E��dk����n?��㬬vn垰�W��m_#	�������K�J�� KʚR#=]v�'d�H./�7@��R�����\��v0��̑V�.�ߍ���u�M	F����'�w�h䴍wRxpYÉ�J��5X�B�;.����&ob	��{f�S5��I˨H�ӫ��@�(S���	��k�&�ԑ�K�CFd*i���;�# ��jr1���J���FO��8#�5MUE6S��1=�Zr+�/=�il��Z��wM���u������a������7�$/�K��t����qm�ٚ���{|�~'��P��*h�r�}
��n_���.u�����^4_��.Z��!꩐�*g�R��4!�ŞP�~���פ�ꃾƂ�ޜ��S=�yTg*!��u�K����8�.�O}���Q���W��{{G<�q��c,_`��n�s�n��Z&8�����I����y����<��p�sqO �R��4����^�׾1 ����`1�o�����,{Wiјrm��J��mX%�Jc�˫>����"�����ɻ������F0�~M�����/��0>O��;9��;ḙ*����Y�j�%�K��3+$�8��P�����S
�+�1����]��}rq�����,��_z���_�{`=�c:%(�\���-jO�o]y^���aZ�U$ڂ��\Y��6��
 �����`�J�0%uC�KcZ�r 5H�ٚ���O��(�S����Ö+��=��':d�L�Y]�"VEߤz�ϩ�C�Õƀ���oҌ,-Im�4Ƽ�����GXΔ�0S�>��ނ���]�4�MThD}k��H�ʠ~FqV���m�69�~ܴDh-c�A!� _��"����5̐�
��f�*%�O�-k����۟0��BEUT"Ϲ�
q�c���N�������}�^�\�㢔��>b��@i�;U�40`�N�w=���R�b��^=�+�#qa��������r閄�G�`]��ښAX�H���Hs>Q�?�O@��i �r�$G��p�~ʁ��q��0{�ͣkGT���-��+�7�:&E$���/����%]tBl��QB��[�Ӡ��s�P�}��
�y���g-I����B�N󞹱z�I��HU<��;�=|"�.���J4�壆��,=�`����!2>���䰣��@�i���e�}y3�z;*�vxfσ��	�`�A�}�Qq��HT�(N�:���J9$]˓�Q/�&��Q�Qϣ�;J��{�9�r��z��jHD��*Wa�X��&�u�ݽn�5��+SR�u��R�VGSB�bWnE���x���d��y�y"}����u�Y�jo��աp�����=�~�.�(#s2}<���>�ATu�M�@$���ϛ9�b	����G;��!^�#��:���t��s��R��Q��5vHx&F*h��,BM���΢���-�5�i��\*�*6�E���~����,tAu��jQ��Si�� ����J����Å��#�����=Kd,��r��7�_) ��e��[!�����`ޣ �EL��lR��J��>�K�z�/�W9GW�T�|�+v&Sg��g��y�d3[b�N�KؑE�x�e�V\�)���b��+@���֕7ʷ, �%!E1jv��'�����4�Uz�iE�^d��Z���k�[��pC��ʵu$9��H�]S˰\�S�D�
%�>͘�������i]N߮����C�N��ں-�u�k��P�/�Y�R�N���L��p���~����!�P�\ ���S���V��r��U� ���2��kk���5գ^�`sǷt	����-���,eߔ{>o��!�5T���t~�<������:�������h��\~��rQYUz���=���-�~(�6�g����g��,j_O�-S�Pߘ��?�d�z5B03?��>������H���(�7�)�x$Ɯx���L /�yt�jKsz��'��*�M�vʻ��z<�cF�p/�9vA���1']��w`<{5To(��k��l�^i��(�[A��cl���vҴ�+%�UVW�7c��"������˸)Η^����$����%�
�ϲ��'���F@H���������t��,K=M��j�5L����)� ,51��i���"����m��1z,!�{��K�`Qh��`u�SV��Y��'~�4�:�-��x�1Rj�})؛�yc[���G�����H��v��M+��_�Aӧs��s���>�u��8Ć2<o�i���u��?��%���[e��L�3���q����5��o��6O��d�ʠ�ѭP�L�O�8ҡXw�����枴Il�!�o��sٚ~��>h�i��?L��0N���ՃX��oQ�W�Yl���^�md8�/��_��6�|��-��?���B�Za���ˇ�w��1���P��N���o�2%�+ܤ��ay$$Ն㕊�벆<̗��ܵ���vp�(CU��g���f�h�W�N�Go�)6s8�#�a,M�ф�Pҳ:���I�Q�����\[5/��?uc�%��(O����^Dπi�5�	9��������}���+g�֒0ֿ�R�E�n���$_���U&��tE���&�t}i}��K�'$SI�;T+��!�p��e���2|�7iD  J҆71��jϰ���h�OE9q�4����*q�����Pͭ�G�ʅ#�f_(��/`M�l���5Ƽ�s��ǰL�Mi�b���d���
9���~y�9M^�g��8���.�k���8�\fg��:OJ�b��Q�2�s�ɵH�/�am̕?@eI���o�-fk��"�I���\�kտiF;Ye`������l.�{=F'�脠��K�8G��s� =�s�P��bD��� ��i�i�l�dʭ�/n�M%F\=;%�M�><�%����1'l�'��n~Zs��5��Y��Q��D��}*���\���ǆ+��2G&�Mҕ�PI�:�^��K�9�Q�|� G�������{�:�u�A}ٕK�L��7��@�f�z���r��>2�݉�ۡ�j�G��n�u�Q�¯����~~赲�@��r3?�fk��7��uQ2œO�V}E�D��8�?j��H3"h�-�Y��d��"7�fY�mN�&�P����Mek����^�ecK�mE�vG�"}�:��S�_5�]��t(�q��Q��ǰA��}�tt�3�s�Z�fL��ʅ��w�^)�>�>��fe�E"L����<p��<ȍ]�Ҿ� �ߣ+ፄB-��I�����:��G��`l�=��3���B�z�����D�x������T}Fn��G~u�b�W�
���f�B�%\j0.]��!���a�# ��e��
�W���G�@�
�W/2O��/!p+Q{�.�k&��Ò��|��
�t��Y���٩MGioWA��7�S6*3�PqO��@���L4�B(�Y �����9�:��e�Ey8_��Bרf�:5S���[[���-{	S�ӰNF�P`HD�Y�[1x2�T�	3�w���p���_����ZҖ�~�>�N�-'�l ��g�㕍j��ׇ�x� ��Y�s#����Z����"���E�z��*B��-��!З��Y��0� �k��P[������[Ţ���A	t�����w�k{L��Y�=�����L�cݔ�T��ysiH�r�G4���GY�A�8��)	]�ҵ�PPfUF��Z�1P�+;�\����XI�]�蚍�N*����b)n��y`�\
_��K���2�n�ȫ���k�̺�G�Ρ`V���'����\�Y.F�4�fn����k�*�+ɨ�)���^+h�<NhH�3�F���OzD��G��q��"����"E�ѕ�r��<'���j�c$���.�3r{c�@��X�jK� EP$@o��y��t��篛�%�J��ĆSܤf:K�RNDc�%�}���߈1���1Yj��%�jf�(�0�JukKm�6��k�Z�|�e��p�ؘ���%CV�KP����GIb�?�0�� �?�?z���Tؒ��T��4�֙\B�<7�ŸH'�؞e"���o���͢(GEp��'�_M�eVz^�b�=<�uXlxVHYEB    5914     f20t�4`���7�V"n��,5{��$"��?*�c6���+�Nƚ$>݃p�]��eC��zv�@�)w
�9m
0X-L��Z�l��㊛���q���5�.a�*�]����>WzJ��n�V�<��{��'k��?�����%��u נe����*߄X�Mk�'�>�߇�b_'�e#�,C/��l���[9D�+�"�bw��@������Z�F�t��'�Zo7j4z�=2W�K5"��h2�7���}�bu�2�Aĕ��[��K��3ðI�Wk�%U8
:�Sa |�/U��-��
��^;^1O_Ch0<��zAPû���L<�5sy0i*��Qa�u�BQ�$O���?�Q������e��Y��e��a�7(O؋!�EFA���7Û�x����s��Q�A_ѰxMS A�����N�Ǯ��^�-)�6uo�4���/���w �|�Gy���[�u���$k�����M>o*��rf��~����d�߀^��2�Lp��Jf���r%��=�LS�PN�f��#%��������-��������{Hb@�gb���n&�y6Ōih(�Ȯ�l��ۿ� o�[	7�z�b�|�M�
��Q�x�`k0�x��r��)O���4��L��R`����
	.�:B!�#B��te�r�.&�G>�yFB���i��$�_�BS��z%�$61���Nt�Ʊ!X�;#Ʀ��I��/ΤOگ�Ս�����%aj���b�ת���F��=[T���	��l����c;�y�d���I5�O�2�6�!�d���Zެ˽�g�>Ú�Z �&�y$c�?�>)������� ��v�Դ��jP���q�K �<u+�GM��ߨ5a4FY�,6Q��c�i��^����@ע�.`��f��mU^�x7��JS}�6�{\F����?�2�?�	mGH f����@: :��Ym>�$w<�^���e��+�qi�0��e������78�����=�ݣ:gy�-tOd��/D��� ��C��F�n}7�U'�ּS���q�%�#ѽfHI�:ȡ�����OG}j��K@�O_tef���и|Q�}�+�7 �^ .����ۨcUc��|kA�DSį{K�	@�om��{���f�:��9BFq92���B���3��Q�u���,
��F%y�d�ݵ�#�O��3dI���1�9��rF�lD��v�LP�q���0%��ez�#�3�o�t����h2Ҩ+�s%�_#�o�r̫Z.�D������*^Y[�g\�=���Fb�ag<�ؐ�h���������-*�%a��[�����	֥_��v��vN^wl�F����r@�=����b.���5ڔNL�/� ���uS�z� �AU�*.��� �Z�D!ŷ۷?���������@��G�߿[���!�iZ���	fÏM�lƖu��cn�:�_�(ફ�go���/�Z���&^!�쑍Ƌ�JT��e��\t:�x���}<Qt�nL�F���xo��=1�x���B=C�-��MC�?SRY��>�����+�s�n]����=CSV\^�<�X��o� e����?~���c+�#{HC7�;�������^Q�0�a؄��f?.U�l�yz�*Ĭ9m6&����TFǭ4��R7�,�g����0���*;�ӂ�,��*[7��I�\Mo��<8���.����ʿ2;WÏ��L_Wv��͚�um���my9��m�(���!���2�6�"�%�������t�x7��8 y��%j3
Dii�Jy!�P�Y3�u~o@61��y�?�i��v\��~�VL�Q�����+�^?�[I֢܊q�;���Ռ���ed}o'�ޛ��[���:v��ZG�+��p��Քg���SO�Mm������"��w?�iPp����4�#��������߳�U�~�ѳ�V}�(��.E��8���c�� Yr�6;+W�c�աR]#^�WMD��������#���՘�]�6�`�Y�Q������f*��pW|�f���h��f�\���%e�6�Ѵ�����u]��Ɩ(�qn(�t�}���I�U7�o�5��o@����E���!��I
Y�C�ף�i��A@��"��If7�K�QaE?N|�l����*���\i��{������Ph I����@1BC.Fjv�-I��A���S�:�e%E���c����=A��"��M��i`1li>��Q�u|���T�O5��y&j��밯�ȯ$&K!���s�C1�+�Vg�Y�»ds�[K�!���"F.`ey�7P򬐱�u���n��DE�ӎ��!.,���$`'�l�3����P�.�&�� \�������	;�x0|�>� G�[ʃ�<�b��
���$�\��MȒ��I�~�K��:���@Cb��C��oX��,	{1�I���[ʋ3��d�G�.@��}�7yW9����|ȦT��ZR�$� Z{�&2��L�֕v.����h�:�u'Qn���6�1B�I*�K��tj��e��6'�c5B.�k1{����� a�'�m�+�v�����1�?��_E��w����`�/UF_;_�/;��H�t&f�����b�HY$2ȹ����r�5��n)��kVD�����!�4E��O�!Ty�v�q#$�Ѷ&1+�q�&��KVL)|A��z�j��\���!�)w�
�TJqZ���ז;��%��a���gRE��ϱ�>R����5_[�z�.�"���1G�<��Δ�/y/��bI�70�U�(vK�b��'v	�z.utK�z|�g���#F�����H��ҬZg5�dD�Η���&�>�oD�,&��8��b���� FI�V<2��$$�6^W�X�|�@�����:���=U�{7kw~H�Q^����y����&�0k�d���k��7�WB}*S_��i��\H����;Ŧۃ��4 ��������� w�!��{9p2�x�O���\�#�cu��!��I0������6*�_�9�3��/To�����x�(���CQHG����x�.r��OM�4U[�@���q?�(�w��W�\�X��کK�'{�\��áI�ß�r}m|�⏣m��S�	䙾 Y�K,���c*)�ȅ���e�9�$
���H�,.�ϱq��ZT��S��8�{Ԗ�ʒ#�����w���q��v���̙�j���c�κ0��.B=�B��HY��$E&p��뢲���m7�s�\�8�$v�ۺA�����mW:.�����s���;*�&��\KB�	��k��y_WٱnAG𛷑D'�Q����H�TdI(������=_ewU$�#ɔ	�%.�f��e�����9Y�@�hD$����� ǣ�;py ��\�ݤ�o��)�m�$)��1W�x	Z��ѽ8r�Ld��箝���^EMPLSr�Щ^4>����z�"���@uRj���+a�ؤr��BK@[�"���w��\�h�fq��;�:�=�"D^	 у�pu��d�I��#�&�?'�9u�W�	�@���?��M�Q ����6W�C ��-�6.Y�=��=�[ɅR$J�������'��P{meq���
ڔ���ƛ3�?�
��`s�xT08Ǹ�q�;�ex`r6�A}��1Th��Λ�ʝ�g�HYڼ6KzQޭ'�T�ܝ�c�����g�*<G��O�{�$��\�W��2<~;��0����C����m�T�JP-��pcv�/4���e[dk��هL�2(�D�_���p�]?gQ�*�1�_&���[x�oB���2�;
�]OK�fv)��?