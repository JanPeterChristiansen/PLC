XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Kq�M�@B(���i��LT���W{������\+�
�bIiF@���@�s��_�}���sc	E�/T>+�dO(�6�ǼyaX��$9�?Ѧ���9�����K$�lۨ9ߺb59c��
O	>h�X��Zg��!��u����(|$�t�_}nҭ+�m�jf�U�]Ǩ8g���)���x}(b��R�L>�@�𹀷�q���txD�J���5N0O�i/�D �k#���u2ݷ���\��X�.��C�E&O���?�gi�\�Ի�ŋQb>یy�Q;TJ���i��8XH�"��Z�{af�,�T����C���e+�9�	3�l�0K��J��E3��`�vES�;~�����^ItN�s:�D�33AI�8y�X(Ǧ��������S3V8Q3���fm��DӲ_����pۻdzĖK�7��6�6		�s�m��h��k��Օx�,���"��B~�{^�F�ןBu��#k�a[�����٭=��Y�7�o]1�ӌ�L[MU�QRQ�9Êm���ls�W��O�;R8��u�T"�0�Cf���a��]R�l/����&��8B���~�X���>�^`��Ch����g��k��bYH�_͏���y>/���Ֆ���|\(U�(�a��+
���HuG���G����y�2po�0c�oa��:v?�)��n���@�e=O���Pޮ�*Q�� =�g�D�F*���L�@�C*黾�����ΰ�z!k��� �qk��,S��9��XlxVHYEB    fa00    2910�Nu��F��+9��?�����\)>}؎Y�L�5�����$C���jb����F�8@�'z΅������PG���?r[,����%��C��#��h']P���<���T3R�2=_{����論D��a��e˾��!u�<C���8G.H�C�{���g^����$SN�3ۏ
�����x?g�~��.-~ۇcg��&j�G��bO�:qBZm�t�C?��#B�Qŗ��8�J��YA�N�[Q��}H+�n�#��䣸���&�*�(]����EX^�p;��������Ȅa(��˪��K�<F��Im�(��O�TMQ��-��:�8ȫw��"��A� ���a� 1A$*Y��@�?̤&�U��̓J4���{�Ml���V�*��`���k'+b��O�# m����0�<	�z�'��љ�p8��;��T(���+�+�=?-ӎ3S�I�q�²���� ����e��p�ϭw�`�������3�b�_&\�|V��;D��E۳	a�A��^�l�U��� ���v~�'RW�����v��?Rty����X��9�K�p��}���y>���Ft�-�^5�ɚpi�^�))=����(
D���5=�����6F(���)�=u�IW\k4�mz*��!ZƜM�\P䫼��G�/�#�j1g��e4@��y�G25g����Jw�rΚ�G�����8-�!6���k�Y�aI����E��oʇ����u��D�^��-�[�ԵN/cV�Y�l�ZR�c�W�s�z���@g%�pg�SFm��Q�׽rσD��w�Y����X>�G�	���)��iTĻQ�?���q& �$	��f氣{�/���9D%�a	�'������bC:j��8�h�! ���}f_�]��?z�&�A6�m;�Ba9}��=ޖ���X�����*��.v�KK��j��`Cuc��J�(��7 R�b�E?�ih�V�����2�W����9��]�J���FI���f�`0
d�y�3q৑4�'�)nW�6QE�5�ހ����9�8U��Ğ��6NHA�5�D������S�]fi;��n��7�/��ғ���U(�Z�R+pX���
�L<=r�������C����x�Hl���J� ���J�<�����f���ao�X����
��+:�D~_��Npy�:���������b��z�`��l�Aq,�j�`:���Y�0�D�A���/F��N�����y�%�
I����\�R��,�F8�&�t�%4�ՃmJ�ҋa�	cn�He���i��J�2��_n��x-�D`R�ڨIc�Ĳ���獛  ܡ�ްoԪ�MB�i~t��D��I4h�D����~h�L���w��)��K��.��{f�U�O7� B~�����X���d��R� ���9>��.�$�֦Ki�ӣc�,�
l�2��`clj�^aja�r~k�Z��5�0�t�-!�i=���-��=��Y@��X�&��D4��kȅE)��!zX��� [�y�K��@�d�
��贌�|�r�����}3{0՗�S�!G��md��(S��;kG��Sdx@�D�<A.r���ŞG8�����2�u�X��
�Ja��GKy-Z��z�G�.s��
���0"5_k���u? ԒB����k�UàPov��F$O(��a����bu�E|�8''��U���&it�D�_�#��}�S�fU>,@ߒ�_9fw����$��t��N�H�J�<� �f<�9�	��,q�ah��`�?m�J\�牢�]r��!*��>�o\O��_ho��G�k�.�b	�x�U�a�?�lK���%��6��n�Yq����6�.dp�M�`_�x�^�����Q��9bn�Ĳ�H��N�Δ	���@&���Im~o2V�9Q�ᘊ�S����>�$`�G��@j�|�{NmH�F ���ϥ�	 A�\����2_�Ͼqs�A�� ��Jcg���R���C��C7h7f���2��`�3`�v��J���_����+{'c3)
Di~��w�x��_[Ǳ�����$���բ��2U�jl�y���4q͓|���7,�t����gd�Fh�uL��*�C{{��p4�Hmy�kx��Dy ��.3��? О� �M4�Z�}/��>.���j�U��)��tƬuwl 	�M��j�p%����~0�T�@��3TH�h�:'e����u�1����t�t��LU��vu���R��-�!4!ȺŐ@��J�|Y&-o����%� �7.~:��˶�Q��[ԥДX�.�)8���O�Ăb��T��9<Z8*R+i 8��9�{.�R�����MY�o͗4�_a���0�uB�a;�Nԇh��K��#��+�w����*�"���`� �Ozs�S+N��1��y��T��B��Șx��T4#�=�ax�"�Q��z����/0�%���J�69t�Ц��e-��b�vd��t�F���_Q��|� �鍦�i�Iq�� �<�p]/&L�~��$w^tw�mW����J�'�M�[����ԩ4|-�\[�7�2a��i�z�v�|m7Hv� �~�]���Űp���o��&o*l~�:�-꺂Ţ��l��N}m�h�A;3m�d��b��%_`����mTn�m�5��/%~V�3��gs�� ��%��p�p��g�B'���}`.�>�8�-f�I:	�:L�<P"dɮN^� VEq^q~�cn��h��^o�!m:_��e=o�Rn�ж�t�V�T&��Zĭ^�hs�U>�D}X���eY��+R�Ү�՚�+��e�#���?F��m��=�*ЄR�M���(�z"��+�^h!/������]L9�?�!�>��`��{�験F�:kP�Ώl�zU���r"�x��F�	�܌��hU&��Ԛ�1����n�J�X�CdOŴץ���2�i`z�/RL�f�#��a�CﾡQE(���C�y�a�����~�M+��"kW���թ�<��YU�sB�׮8�)��\��V�6���a[�˒D�I��*ު�w�B�	����W{���8�3b/$)�M5�5Թ<�[�ʮ���ftrj��(��� V�~2�a��u�1r2��Y�%��%�n��5՛�U07�:��z�o��M�)`�c� [v���vA]Uyս�1hx\P�U"�#�h����G���Ѵ��8�ϐR� =H lx塷�K�6�]��3.ל �nx ��� ��!�������T�|_߳
����'�8�n�-g& ���M��%��tsJx���sl�f�[�	�p�v�����.�G%��m}������f7�| Y��n���Ǳ��3�2��y深�ɉ�0:wȱV��@s��Nd�4�@h�>w�2�|5�͘ ���O���<�Vۘ�c��C�����aL������Pꮡ�~���'��³p�{⃶9�5��ITE�6A�y�|��DT�?��Gܶ�Nt���Y�t߲���gM���e*p�΅��x�9��9+< \Cw
mˌtA�v��53����n�ͧy�C@7]��G��> H��[+������'6�OP��f�x����/t	.�>��&�4�~�n��Z$����)�D�׼�5�R�H��k�A�V��m��ьK�*�|�3��������fϩC��_��,`v\����|�0�l�|��k��/:o�uin�#+B�P]ܔg<��_g_�
��~�S^k:��(9ǝ�ŜMa�b��으(�8u�R�`�=��Q��I�>�[��HQ��n�
���e̜���j�w9p@�H�-�C_O�Ǔf�]����Rnǽ'Sӷ�2��c	���?�ڹd��B��&2eKI] �=��#C�{�ǣ�x�j7+Q����oU8*���#{��_2�������O=⑦;ҝ�^�Ä��q�om6-�L�c�������@Э����y5>�"����{�&�����CjH��թy��bͽ�=��*l�\��x͂���+1H.�bE�~�魄������F����ceH��ϱ!h)VY��1�}��TϷ"�X.&�E�(�y�t2�L���(Y���w,]��$���B�L�Z�Ɨ3�̂|/���x^p�a1���M�����ۛѡ<���	ՠ�a�gV�d4�§��R���Z�S�}OfO��lƺ}��7��/�Wj՞g��m�5}�}2��t�'*�Q�M߇MF�j���f�m]~�Z��f��0��M��\����kK�)Ѿm�j��#m�/�}u���ٱ�c�8���g)-�ḏ�Ĭt��?�"�J>�ᜀ�}?B�M� ��F���ؼ�$vu��u�7p� b%�g�����5ȏ�z~�$�^��J�H�$"�l�z�
�~�[3�|�5�Yj�uNo��5R�n�8;�̠7Q��"\�Z�xQ��4v���t��o��G��������(s��a�ԗ���	�]l�-z
�^��ʰe��u�ڮg��Q�ƆS��蜰��,��MF�����w�2D���(L.fm�Ѵ~������ذ�?�hB���0��
dYw̶�l��.餲���i��-�e{h�Z�М[�n�����3���K��ĝo���}��?�_��!*+f��141����4<b�}������dd�ڈcR5�N�/=��mC�N��N!�:){������F���v�#�Y�F�l�e���k��l}*�ܑ���ۂ�d?�a���=��`.嶇��V����O�����"Ԏ����_�NVQ�T�����ED��^���95��k�V��C(���&'��-�����Ŏj�6�.Aچ=<~4���������L�8`�A4FA��b��=E�)�$�OFKx��q����My����	�6W����
����Fe#��5Nh�qߘB	��/J"X�8����ϸ�N���(��'�A�!C�g����r���XK]"Gڇ7������/��r
���"c���٦�@�ٌ�Co�9s�{�J��'�{K���uKY��vʴ���7,��k%��nU�|["4ʣ�V� ����abѩ�
h�&�8=��%�ZY�7��k1�0����k,kGR8�XOq��;���7Sc�q�}>6���v���i��K�
��Q'��/�*r��U�5 ���5!f;N�k]�C�{���*��U���X�z�"�n�m���(R[f�H�K�4*��v��kl��-9����Q�z���p{h�O>��Z��5�Dk(��Dz��f���]��Q=%�l	���m��n�oi�Ő
��M�Sy�aO!/
�3���U�z����'[������=k	�m�}���s�ѭ/�i�� (�8��̐�E�%���RvŖ+F�>'E��veM�[�����m"��ˑmR�[�Mp�/ G����V'E2�;����cA���/M/y��j���m��f�Χ�Q����F�9W��1�W�ƌj5w�xHpV��ݵS ��(ߘۢ��Β��ap�IS�C�ڄ�u��7<�$b��t�s�lc���L<����1�L�3�2cyZ�~�L/T��Ol�x��]��/�s���$�����tf�G���k��M��!�IEݙ���"���h#��(xe��ˬAfU��@��6��p�����2��b�����1�_��WKf�����1�����q�3�uN-�m�8��/������nٿ�R�=�%m`���Ǜ�B���Ċ�z�p�A�Ƭ6����I�"���~=)*��Pt���+�f@W���p`1�*pS�~����O�@BO���Q5$���jo����<�9�x#7���Z�z w43W�OC��w��=��'g�
̲{�Du��W�ʙN�-�5'��W����n�z�y�
�yH�Bp1�=~�u�	 �ˆ�̹u��i"$�S�A����@r?'� �4rd�b�p�Y���N,��F���}�s¹�z#L��\�A���4<CmD��okh��U�����z��h�ҪI�Yn��I�v�_�Ǟ��� ��F(��c�b�%���W�	7*���|м�"���'}�ȼ�
�UGN{��+��/�]Vf��e�!�C��b�T��0-Fh���5v�]M�216-�RM�;�h���r��k��
�kn�9�����2�!_�%���,�p�6���	����E��z_󝠭%���M�W+E4�Rل�Cz�g�۔{�C��q����Of�Lw���[��Y��{���C�i�s�3݆X^�������2�݂O�Z�v��7��/�5���(��'�!�O���_���ʏ�Y�)��;��}��o{�Xy�<���Ҹ86��D�&�V������k����dې{�ﯹUVi^XY��l
�ȼ�8�8z����f���/z��MX�ٓ�j\q��F��������T�]?~���$��.�{-�W,�t4.����� /zOw��u�n#$
-JjcR�:J�#*�t�o|)��Rz�Kϣ�ծj�Ÿu�H͊�Qr4�y}�C\H��s`&��}5>�Ǜ�!0�2@p����)�8s������l��n�_�}�z�9�:�T�n2�+G;o!	|��TV��hx�r���nn��]T���>e�T���m�8zz�ܡ�~�tbI���B>��sFE����<�򪩐{/��)4ځ����H�dHE�>��<����9/7���;�J3�[<��$�M��a��*��ꩾ�Q�������,R��^���HO����l�7�G릓oF�1���̋��?��:i �mذn���u��@_M��LF�	�(��K����M�_�<��)�Tj0�S$&�A!V��@��2�b�=���~[t�K�t��G��������@�qyU�uT5�8x����ټN<Y���?2;��� �>�R�YI)4�d�^�*�;��;[�S�����M�D8��]�?{��#�V����$�j�&(���K�F3?|9���Q8V�9ֈ
�!��=�QT�eGe��U*]	���'G`�]�ƽ��)-D�(�x\����jJ��>%���=�lpB�#>']�D^/x�#4R��~��?FĐ�G��Vhx�)�K<ŧ� ��A��z��GOR���hPM&I܍,-������o�!9S���}*��9O�\2�b*�i�Ҕ±������"E�<8팞�UF�Ꜭ���I�Z]b�n�&��ڈY���Ұ�p����qפ>˓Tij��R|/P���a34�;��ffz�)�W3��1k@��V�L"�+3؆%`ȉe/�w# zܜ �/�{"u0��Ʀ��h�0�9�����o`���ҍ�!�I������X@ <�d��ۣ�@��ҩx��⟬��=x|��Uɩ�5j�ĩӣ�')��j��L�=޹yj����"��;���T�m^Xb�G2?R�{�g`��t܄ųy��ug%ߐ���?��~�K������2�=�x_�Whj�`Y\�#��F�+��+6��a��*��u�͠<��/~M��^�t���+�b&��s�Fz0�V㣦��=o:х�[�c���B�Re�X]�V���/�H��?M���t��!����hè�V�W��Jgl���9X�a�7�}�ެqi2��b/����a�M��������P�~Tv2舶ˣ��6�Y��x���~�y��]a�U���s�>�2�o�A,>����#30�e|u�U �}�Lk���j5�\pv�R֜��ĸ%n��s\�c'��W2ȕҩ�S!j�����sT�4N��\I"l]L�C�d@/��gS?���jG�5aŰ9d��՛��hQM�6E���Q�t_���U��^I�-w��d㠙�g�r���jt�]���
t�O�x���w\hmr'��ŪE����9���P��r:B�FaX��L��Nπ��h��C�黹�6رXP��u��S2]Y�L4��;�ӎu�0�Џ_���S�g�|G)��!Az'�/���HҨ1��h�V#�Ҡh�������x,�B���7�do��S��2�/�v0�`��l��j�raU>�e�"�����a?m�F
j1���ɦv�!'My��4��p�r�NÑ3�@0M��[%���I���c���c���mIryIP�Z�D!%�����&|���
�5�E]�ە�7�DZ���!O���g�4�3S�VO-�!���b����p�!8��?����y۪C�縆0Y�~fF��b2�����ՒT�mY�*����m���nT�Հ�"�-��@(����WK��ʵFׄ�e:Kߴ��A�ǥ�h���{Ͱ��>ۏ����z
(��m��$"���S�u�~~�t�6���R�����J:q���)�6��%Xy��H���"��;��r֦r�dX�8��V��f�di�WC��k�%d����Jd59��5<��N�|P���Wst� N�^s���j%F��H{<�`�>� ��D=�����Y�W4"ߥ",g'�5v.�;����c�e:-��p1T������_��n��~G��=.���Q��7Gr�ރ�������?�yy,A��������\M}n�h6L)Z��7=�)��
Hp�Y��Hq��el�\���"᩸y�}��1#b�i0���D�˹�TW���H��y�X�h����������r�/筧�NI�w'	\��ǝ�Q@k�~2*����k��?�k7uy2�9iM��HáF\B.|��W%�[�W:�J�r>-�D�������Ly()�?�x��t%F7Ά�y��d*!'(�5�rgq���q>�Z�����j��BB7���"�≔�M!/m�U����(��e&�}���	�?Շ���j�	3(:�f���K�;��RH~T��4����g��^�m�5����+�ʃ1
����qh��� �u�aDs��vg��qJ'�:ƻ���8��Zk������JB#d����X�az��o�9�s_R p��a�5�lma����f@ژ޵1`���5�]҉D��3����OBG�T.D�e��W���ʶCH�m̭Po�#M������rT3i����a� ]g�rB��/"�2;�ȟ��lQ��� {r%Fyk!�J���g�ƣl�i��gv攻&l<�������Ăe��S�,��!{�e�i��Qa���!6���̀?_�ډ0(�����c�t^^����"�s>�X>�75�� Z���ۄ����0E�c�k5��)���v�d�8'�ah|�7ڔ�^���^�d�B#P�ө��M��}
�1vػ0���A��L�P�H9G5�D�?k�Y678�u���Ӕ���h��F�M�!��ap���r�� w��l��W@ߩ�2��_�SX5�b�S�5���?T�XZ�i��U~5�7%�|�WC�	�О��R���q{�:oTA@CD��>���4@Y9��X���ܚ���
m]��y���Ъ��H{�7I��w2�DNz.!ւ]ܐ�~r�eL��`s��=�+c�|P!W��M��,��ո ��4$󻘥H�����<EW������&Cb�P��Y@��G<��:A��	�E�z����J$�Y��=Rps)�C�:�j1�~{�;i��>���ud�_���<�63���a��f������,(d̸�g�%���M�:�
m����8��*r����!j��c���T����pFAz;�8��V��'W�\�gL��y����I�{�i�C �%i �0���=((� ̰l7	��&�X���C����1V�x\q�N������ ά�Z59��$�ߩ?�hR�:�t]J�ׄ�j���W4��� �U�*��/ԞMUq��]����#�	X���$�[�����\!���R$�&��T�j��pT>RR!U��w�H��K`�Wyf\�l7��4�M�%�^>�Y�4����EL���E.��q�>$�<8�Y��24����X�2m��l��D>����j�qk&�NK�,/��lڥ}�O?2��Nt�TeʸE�G>q䴷*N�	�'jrı����7�0�]1#d��J.��y=��Y9�{�/�SH�YGެ������'��n�d��X�!C���IM�~���ll��B%��՞��LYMZ	7U���J��8��
@ �fei�=�
�m�|����7E���si=Y�h��1�Jc1w7/�Nl��4�`Ke
�(�Z�-��m���B��t ��1���t���Y��v[_[jD�����o~���XƃfT���h@S�~��>#O��3�bʸ��-p9��܁��
��6*Y-npɮ܌56$-f�/S���vz<��]���j�֑O&�ɜ6{8�mX�1�����MR��XlxVHYEB    6184     f80�B��O��PN&O�R_�@4�[����׆؆�i���vVG@���T&���֌{ܟ�e7ƪ�<����JL���t�M�C���q�~����ٲH���:'ևk��Rs�l��OO0X7�ɨ��K�G��j�����6c���M��j�-ǎ���]�=�K�=���菣�� PEꅶ]�͏V9�I�՛l��)��ˡ���v/MEr�|�:�!��G����~N�Φޟ�a�5�E� ���y
�L��S�HEG��מ��ewKr+������#^[���3�V�����f=l�$ �y{���Ì����c�����%�̛�Ml+��������d��|����c�d�����}*����#��^�f�K�������(�y��D�?@g���RBL8$�^�_k��C)����+l���|\M�j�E,�y
�,k�M�|�����gĊS���w�q?�M&�c�2��1���������p+�ZYfj;�@:��&��{�G���m`�*���%.���E/V�.�&E����o���~Ȗ��H˿�r�>�3��4��h��M,��3R@���_��L�>�)�Zے��&٦�$YU� .yj�7�QW��ņ��z)�h�-��S�-�����yTMK���Y���|r ���Q�@�׫��>��4�D���XvY��=]q�x:9�b���4:k�"���6�u��-��s3�R�n�9qZv��̊dR�tͯj��`��]�xN/<��|r'p�8Ǡ�zE(�ȖWhݲݖ�#������`��qQ�lԸ�
�#9���w`���~������_�,Y�9�T��m	�P���j(�$޹�4�}f��'�n�&hB4!�F6�w���xz��nt�;��FH�]��ֲmC�_�W�	�#�%�d�<-�*�A�h{g2�[�~���ֲ57�љ�o�9ױ�?C���|1�>9-	��tŉ�c�̘Ã�R�!��҃�/;8�r]m#[�RK���+m�k�11U���\:��T���p@�k��S3�Ɂ����˱1Չ*/lb�v{�!�4�3�B�e��H�=5���s_!ꩍ��J��V���$��^��0�N�.�M�-��N�����#@B�o�}C{a0+�ʽ���<�O�
1��0{y�C��XO�[���T=��c�1諝�.OR�_��J�/=�AH��O�؂0����A��	ڽ�N���Gl�&�@
W��(A
�@��T��	�wE��<j�"oD�W��E��Ѓc��'��b�y���	L5�[uF�'h�j#$}����W��ȍ�{�7�� �ԡ6��ꣅ�R���oOi�n�(Sz�����^�%�
��U����.���P�[C!wu\������֔�>I��^�;�m5n����H����}�y�#����3�}�J|�_0�G��ox&]�9I8ICŋ��(D���I�%�=��\J%��]��z���̲D��p:A���[��4�l?�z9�W�[��.����_y�����'cď#H�s���w�L+u�&W��u�x�	e^����k�yDtR���2��EE.g	�E\DҐ���R�.��^�)ҝL�s������������9��$<��F_Xt�5��29��[�.�A�)�hk�mO���*�ݸ�@��a������ ()�

H����ii�'O�{(ԙ���揥M��{P�*�<A�����|�£�p�d3�݉:�7��g����אv����[h{4�.�� Wtg\7<��X�WA�-/Ɂ����u|�n34ڲY6�Cn�����jR�̫���H� �n�?�>k]�X����K�T
`�������Tm���B�Pm���R5�����4G���ٕ�xs����m-�9�K"t6&�)���w��V�s<X�ͻ�i� �_]��i>��Z������g�� p�h�
��(d��$݉��;tU=*9�:�q���W;bU?�8�����&;r�I��"�6��Փ��¹�����ιz�1��wrp!D��X�Y��?�#�&P�i�	t��uG�~�ոw�ժ�����\���A�9���t�H*NΥ�Mm��9�o����rY����QL��+V���c�O>Q}"�Bd���~«��PD�ǖ9B��z�<O�t��Y� �/�3�OXr_�gK��+�G(+��#;� >�$�����6�V�+�� 39��N�24�)�?N�y�y
������h����T˵��F����x��Ad�1�
!�D�C��:E?�Ox�h��4�}4�~���Q|G)�������Y<��@�K~rЕ�����̂��T�jۑ|�i|�U�Q���;~I�tb�әd��fڄ8�����E��o��
����9�@^ޚ�� ǁ�#�sS���i�0�pS�k�#�sycz_L��/"۝XZǓJ|�.��9�	����y}��S��`��5S���2 �ܖ�xƸ��1h`��`Cy�;z8�����w�:��~a:0��w����k�$!��㾏Z���,
Ww�^U���c|�U;��圲:|Ykmz(Wˡ�@�v�d���u��g��@!ݲ��a����f��0A�g�HA�a�U_�?��B�I>���[���P�8��lg~T\'���l�j/hY���U��H ��a����u�lfJ{֕4�I��~$i��ʴZ����iRu?�-��D� �	6)|w:�U1�,�;o�_����&���^ �r�Δ���$�������I��P�2-D7��y����C8��8.��H%��_�*#Qj�M$%ʡF�}}t#?q�o�ΝV"Q��WpO@[���n[T��V�nB�[PC���K=�R��7��Lr�~��Gf��-��vІe�i�hE��If�\�q ��e�`)�<W�=�նި� �m�l`Vo��0<���l��{η�����"+#��H�
=D����.���ǫ;�U�Z�T1���v�3�M�7P���	.�N:�%���j�WVc�����F�}W2`s�����e�j�02��b��QS��p�NZ���c�Ũ�xJ��qa�A�/@y���fog�uCq	V\�W��܏t/�Խ緬�U,�*��-Z�-��/i��}�[n=��;���&�ߟQ���N���ۢ��Պ�*H�uP�^`C�?�F��Cc���Y���6�s�,
h��ٹ!����ƙ�Ҟ�bɹ����n�$4�u�����R���I���N�)�J��� P�L�y/�d��b�4��I��ٟԉ�=�J&��w��A*
��)5�-���MH��r���-u��G��=B{�S^��2��۱��H2Q8�iC�M�AH��-xIF&��� �Q��9�c���q�N�Ǆ���qDx��܇�G�o��΋F��~�K*ll�rvi%j��L����5E%�c���p�ŗ�<�h�/L�z�L!J����q$�U���al���Yg��#|�Q���n�]\�ԌJ4.N��|r6,g�@��"(I�rP�Ə<ƎuIMC�jk'9�芥��۲�IK�1�*(h�K�ե�Ad�x�?�5_mAX��n��L�!�p,�S"��ǵ�@C�s�v�'�ǟ����R�!�T��y���%�f����=�%���	g�5-�Z�BRs
���/1�g�?
:�ei�;#�(�}������k�������	�)= ;����3�+��`���MV�G�|���ɖ;���sM�����M5���-vˎ��Տ��w1
�]��R&�$c��wʴ���D"���P+�S�5��\|�L#�tK��]�m�9<��hqI.����<{��3��C�����X�J�/mв�C^x7k{���֢D�w{���E4�!�
��#pX���銓[�I+K�dGI�P����6��