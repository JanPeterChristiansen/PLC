XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��%kŠn���^Y�\o�v������w�j6��I�{�� P51�w�䁊�H���MP���>n3�6f�\M8����iQ?���gSOA�O�T�S_���C	�D���(ޏ�'"������n���[�'+��*ߔvO��M��|Vis� �ω�ﭡU�^i�z�p�>��N���r���l2����Y q��,�K8�6$u���Ŧ6=�BW�:��ut��K��M� �aj��p�A\�nR*���l]�R@��X���`��*b-* >�o���G��`��Blc��0��6nl3���x/ 3���+|u&b� �)G��V����,b�6��{Z����P-�π�����Zr����JW֩>�A�yGS�[\�%*c���R���dv}Xkg����̲L�A��U� �S��C�M����y�	e�硓�$�IL���G��PnV�������v�Y�|���-Ñy2)��� �}�� ����]Y�:䲨x���X��1�*2ЦnD�R��4��?��ru !����C�EHt��W{qj��HTaX����b�����3��$-l�Gk#�rZ�D���l�,X���1a�YH�y���_D�Qh�%k4��aR5���-(n�Ţ?*o��S+�n�\v}n@r*>���Vf�'�ׂ$�Ñ{�<���+ C�� î؛Ν�ϸ7�؎�/���R�г�����>�_T@"R&���_�'}a����L`l�`1�'�ɦXlxVHYEB    ea93    1880��8k���G���r�Nܲյ(����A��E�W%=eCEk�,�X���1����A�sj���)*P�� ��X�*�"X-^�g���-���A%r �X�Eڗ�r�����c�Ao*N&���e�-4\�EBhYLU�r�|V�I:$�.xԾ��%��A�����Apu��}4����G۝Uc�<�^aU�C�(	Q��Uj
r��jãK�nN�c���fJ𴞓�j��D ���D@�������\Z�qr' M��7@�q��<,����>�9d��J�Ͽo[A�.zT/Vw �xX(0�+��L��,d�êx�|f�EJ?ˎ�_�&���$���¶׀�I�[�بBd�i�pR�jt��s�랓��:����D�%�����*%�Х�^]�#6�����[.UJ2�dq!��>�E����*xl������8�*(i�dC��<K{�bTϕ'!�O���[��pZx�+��"bP�-����d�Sʧ�4T�.Y*D}�a�%s�B�[�Y��@b�1�� �"]�J���c'�K����3Cc�> 쏇�$���z�*p���~�����P2*��V�Q��s>��ԋ��s��w7��3��*d��FEJ��,��Ec���>���&�j���bkU`0|�S(h��=3�]a��2v��[^{�3\/9])N좘'T�u����N:�c�JyŐ���Dh�=y�XF��+fq� }���S�v��.ƣ��dC���,���N�%
s��)ЀT�
�]�GLqz�u��m��e�z�3�z��so&�_L|�oN�x���g��S\����r2d)e/>i������n1)�^ʁ�ރH��Tdt�1��m
/<Ŵ-U�k`�=$�-P�Y������%h[�o��/ܦx��5�kSP�7<#plc��f��iH�x�nT)�*ì�^~�
��dNx?j	��~���Ɗ��,�km��=ulm�J��E*���n�֊|�"|6�Ev��^���9�l�X9�+�i�[��%�1�5ۺ	` A��iXLF��D���[L��n"��D ���	��\G�p�����4$8`��S3��e�)�Gm��v�_̥pP�VR�-cA�
2�UM��#����[��'n��]Ц�wA��$ ����C��Q�F�C*��Y(�Eďx*p�o��2Eo�m66���ؚ�Ñ�5'�q� �0j����k�������@s��+/�g�ї�/x"[%��쒯[������x f�[��v�̞�����0�Ԋ<9,\���4ڝ�*�7��|8���ԣ`:��U�ܻ�?��´����EP���Δh��IP?~lz 5����I���'+k`��/�f=�:�t9G1�JK8��Oui�1g)ԉO l�? 獚��S'?����ڄ�D��:m�q�1:N�7&�T��k$�DZ&�+�R�F�|�侕��S�y��t�{x��
���x� x��O�*E�e��9y��UUP�����4��]�|b
k�s���n@�jW�e7ڃ���)�=���+���3pwū/}�AsBb]{��(��)4n� `��3�h1�­�A�K��-����.dM����vr��"&���R�:ʫ��J�|Ιy������;_�g�H3|y�l���$���-Z6ṁ��E��]>�!usѤʠ-�5���A��"t����c�Y؆o��j�6���gY>���vH,ݪ�ؗS�D��2���N��:�XM<�b�L�*�k[W��nh�[V�>�(��ZA5��iE}Ɲ�d"~���@�"���D~��qN�|W���).�Bnx��o� [��g��)���?�_^�����\ş���n���nS�svְ=�@k��@�O�קF/1�8�
�չ������b��+��`�a[&v]�띀~Abk'���f�=.�,P��.�U�3���!�?�C�.��;_l����HC�(�G�Ǒ�F\-<Y'�/����̉&�0�X�Y�0�j�˙��<�G:�[�Z47Q���f7n!��q\�>�5�K�<N	����?�<
�RC\�Ǽ����v�܃�y�Q)�G�1y(j7Eb��a��C�%��}�輫��(~Y�|�PJ`�ç�F�����}����JTz%����9e����Q8+���f�+	���P�*_�DGtS��׳Ē��ʒ6jQ��^|�
�>�v��k�K� ����p2�ll���nN&k<&��ۘ\ H��tU����Bi��EP��l!�[���O	9M�&���7����ʱ�B��58>�.F���~A�I�j�ITy�_k�a�Y­�@^z��mB�痢��������Xz�9�9��AlO�L��3и�2��6f��pO�W�҄���"xԀ$�k�T9Z4v�/)� ���2�7�͹�HWm��x�S*�F�hZ����"��|��zj��[�V[�ݢF0���"_zS���ވ�B~�ճ-���W�!2b�+{w����,�!B��3��uj�0 ���lK\�p۔)��c�cj Jפ�7�[��N�ڵ�L���^rzg�]zc��J�Y�N��m����o����#�G,tI����6��_�/���d%��� ����&�~m��JX18���|M��d�Ũ�8\�������_��6L�y`��0moLx�;੨k���x52I�\�Um�����r�y��mSsF�8n~�D�rJ.u�̪��c|/HR�{�{ؖQ�,�E�9��:-��Mg}n���O����m����a$��!����j��:�a�Af���d� ��6�uǶ�O��/���L�&<#��4�P^��Xz��2`��A�=�_�c�~��&�~<K�����ߤz;��.�TGl�4�64���]�/��������X��m�\ݻ�a��,�����6�s{����F7�`.�ò�P���o��H<<��D ׾cL)_|����ǻ�<�`0�n:EH���B��u,��h��얡�W�DL��ʴ�%�؏\PA�<�{D�	�����$~�R�9��S���Nݠ?	�|0�/�7�_t{���؄�[��t��*�g�+���O	�/0�qM��ǂ��[��n�*h�8�M��׾+��'�6W�(ؐ3���Ѩ#ȟ�v������~1���A-���x�}Q��`�ݖ�D9�h/�TShgt��~d,�z�����k$�z���q�X{��#h����N#29l��D�~��lb�҇s��0�1���e��_س[�Z+MT���a�p�1��t����|����0c[����p���o��n��'[�b����y�1�.2;�v�5e�N�`
k�=��G�%�]���ݨ�?A¦ψ3]��^Ky��]1a�����1�íh�����ꐲ��d[=v ɔ,�n�	��"ve+��I���l�y���Q�`0����ռ)�?��PM+�^Vg9AC$o]�D��i��f߀A�@��"x���=N<}�`g��0��G�|����y�fs��^뚣�24��3����
�d����y�:X~�k�����$y�H��"]�s�ov���umI�����k��a��v�Vs�N��4�� ����b4Y�~�kQ�<Z�em��uۺ�SE�mv�Ȃc���?x&]k�ꔚҢ�CV�2LU�Ih�O����{7�PkW\���NA�6jMD���.K���-�\82���+�#[E����&�<�RS��~���}
�.2�}�4fnOZj�|R$�)�c�]��Tnd��z��9���"�Bg�*6gӲs�9�XU��{�C�Ә5���>�����mu��C-�$8�����x>�����ϛ��&���M*	h�"�~���9�}S?�ġ��uz2?,�6$���� 
�.n���6�0�S�d�>�]bm�?�wO6c�z�]�c�Pa)`�i�y�E���āHˢC̚^�փR7���,��h�F���Gh\zR��%FT�&7%j0`f���d������
w�Mi�����˿Q��{k[HG�eq��0T+qfr=1�S��V�v�wmr��^�4D1�9�����c��,ȝ�`�;����_���=�h#{���e�K�c����N��Z�8Bj�|}��Y� O���LP*������sE�z�Lں�!E���%�90�Q0U���,a�h���l���ǫB�z���S'�!�c��l��!-:���_�~}���1��`a�� ���[��=ש��ސ����G<[+�9w�,�n�[v����F���1=:p+2���d�D���t=`��,ޑ �)&��UqV���䮥ĩ�ȍ���S���˶�
j؋{�Çl�*�
!680䥌R)����8���pkj�0�w_��� �:�ң��m�!$:M��Ʃ��n�[��]{s!��1:�C������O�d�t�	Z5a��_���M��|~��O�Y���S��]h�W�� ��3ϱhu�|y�	��To��&�4��FAb�F��P��/���d3	N���Ds�������֩~�om��N�?���0F� �� %[�"!vK�Eޕ#�e	,�N,"��b��H��uZ�3��T��K1w�~����;��΢Q�C�Pv�V)��ع���G�׷1C/�5:8s���E�鎉�L��,��g�\M\�� ��8���v�9�&��lՠ' X��	r����g���e�$����՞��{	�,���5�����@\��n��� �z��3/�D|`��P��9Ъ\.�y@��`��@~HGP��¡sW�69��3�R̲�(��W�l^���8�1T7��5ͨkC6e�+��5�p��	�q`��]���_�;8��w��Q�dD>k_�: `}_�4ؤ�1�d�b����K5"Ty!��u ��߼�k՟y���Z9
T�I
��+L��;���\��q ���1�m��L��D�+���󖪓j�~ d8�6@�vJ��k8�xY"ji}.+�*���r+��hT��+i ����B[O���F#�F1S&��
nHoq?�'�l��u$z�^�9|��8����?����ը�ztz��6~|[�^�������ΎH(Y{�˾�f��ϋ�)#�ƎH+)����D�,#�z����x{_Z��>+\�Jb��Z��/���ά8Q|��mh�i0�^���~�:i��b�O��� !���"X�>���^h�X饾�&4I�s2�T��\vNߢ�?�ǲ�Y�G��☗� ����$q�tۙ�����m�k?����s���
Qi�'�[�M��ޭ���z]){�6����z�q���&ŏ1����V�����M����YV�}n��(S���a+�j�S�NB�^Pn{��^[��c�B�+���)�/���(�3B�9ND�V��͠���8Y�J��0b�7���+��N��~�C$�մ�A���� ����������o�0
Y��I��צu�Shz�r��P긗�J4f		���:0�2ý핶�.��� ��<��8~`n{_��3����z��N��rM��BSS�k� b�*�{���!	�b��ޘ�S�=Q	`����Ɂ�f�s���wY��Yg�LZfT_Dp�c�Ѿ���ɀ�L�sk��FR�.yޏN��<۲P�Ľ�n��F`�B�D��i֭2�Ax��������1"�v,�>�q\b����̷rJ�!K�;���ݯh�K����+kj
bW�{���-�n:��hh-�	��b�G��#�.   ��jBq��]���p"y�����2���}�:�vd�/��S��[v�U��E%�{g*�P9)�g��
N�1��� `�9�7��({r�{/d�T����$��Q������qC��:�60�IZ������B�x���m��q#��r^����:F���w�/�Vj��შ@y^�*��ϟ��7DG~�w�����r"į�1cJu����\�m�М,�3��;0�d@�B�E��O-�\�����_��^	����vB�H�� ���p�k���Z�"��S6�y���Z��n����v���#���Ϧ3�/&^��5�(|���L6�*QrqI�{��~�т�):�Pvj1�pR�l��]mc6��j��ʊE�����c��f�<��=�W!z�%��FJB�����F��?�.�w�gԂ�)~