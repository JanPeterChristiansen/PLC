XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��9����⽆�y��pl��K1"��TgQz� u�Θ��n��x'h��j[}������k�X�f�����Eظ! 6�H4��Z�4��k�L&'��wD�d�����(��@ɞY��(���
�7���M��ou�͓4���И�N"o�F��V�X[��nc���6�S����s?HwX0�.��H�v�^��,V�PO���BH-�|�Kv>�r�1�1��A*aN����ߡ����6z��ز.`��q����اM��DV1;��H���ч�V���M���1}r��un�_i��\�j,YZBw�<��U�W!���[��g�+.hEu1e�'�ɡ'���7?�=-���d#Ri���@\��T� �zN�aP���){�_��ě�����&eqLA \w�IG]ƟB��$�u�c�obƁ���kW�����;yי�4߱��X9z��Σ�!qI��L0ͅH<��t�>��u"�;ػ����zg�:�@L)!W�Z*�Wl�0Rl���I�y��\%�]�P��
�Q&Q�h��&�T{�;��r�Q
����lŗ���lDLeJ~�0�� X�,�Wi*�G����C[=�p��,/v�v"��T�n�:.��<��h;�a�����s3)ܻ*��c"E{~.T.x���:Y���V�$0��;Y�W�97�g����c٬T�=�WC�	9�{	�I"�ȴ_��̶����j��* ����9�U���Q<a��{t�Ε	�׮Q.�XlxVHYEB    9732    14d0��50���v�PdZ�����JQ������׸�'��!������N�Y2��,x��A<��g���X�F��np���2�/.ojzct �	0b4��_K�]	*��܁|/��v�/�X��%'#Hr#<���d7������-����`���1�-�7�Y�h��B;2G�6cW �G�bL(���z��%-'�	��)
"���^!7��&�o��������C{�VX����]���	m�i�/�Wj�ӥ�,?������I)&�'���nc��Nb?!�SY>�t���^�nI�p!Z�Ha�3�C&�����e�2�5��*���$���~�M٢`�9� �TtP)@`���[י��<l�?Y�]+��n�\�
��h�nd��x���~����S ��9�V,��#�(m�l��4�14q�����aA0� ���#��'7�yF!��A2-��"��n;aZ�s�=B"q&u�<�+���N�x|��-xi�VO�Lp�����#\�|
h^����kKH�������q�k��Vv�r�KS6wj��e��3̕�6o��֝@4�c�x���ٴJ8�A���V��:�W�1H'���;�OƄ#��a	����i.����H�n��}P���(���gg0��V�Q�
���R�	%z�Wy o_��%���:!����i�5�����VC���,�j���-(a�4�,�%�޵a�)��^b���W�k\A���	z� ��"�?�Q�G���R�tz/�!�P�ZzB�Gi�56Q3�|�-�o�ޤ�v��54�!e-P�%���O��/��z��a��8'sԹ �hS\}]hJn`@��f���3SZ����@��\�TLR&���G�UUvy1ǽ��~�uJ���y�z�\�Wy�eU]��	}^�[�>J��C�ű'��ߒ,P�;#��'"GOJ�~�����<S����f$�|4}���W�Ÿ�E��/�I��`޲c���ȴ���3�iK��F��=a�E?�����i)Y{�Q7&S���?�e���`�O	ՁY�U�H�K�g��<A^�5[����΃Wܚ;�X�+�6����c��HK��)���'���j��,���/ă+`8�$ᛃ����o�]%&�1*�c�����p6�T��屦
�X�/�e$�0�;n�A�.�ĳ�����ߴ�i^��Q��yG�!������3���t��7������Z��R�����m��i�%��<5����x��f�Ү��Qv_�r��Lj�Pu�s��q1���9b,�]%{s���ŷVؗ%y�}�����6��V��Lz�-H�<�`pO���e1;a?iCx%
p �i�Q�}@D�'� �'�?y/=�����nmV)��OF�L��1v=d��Dx�U�T��֎Q9̐P��P�9���"��/ڮ�� p`6�1�s��U·��[�qy�jS������+$��ĥW#��[�m�Ax���ڮ��?Rr���gSx���Vm���U�߭:$�������&�Q9y�Ow��x#���{�'p<S��U�9�56͆�T�00i<W~��ѤxxڐU�3>@���|�D��O�o�N��It��/�ܡ݊YZgʁ�(!;7;�s�T�,:�����=}�+8���2��/y#v�h�2�����^<,B�8�V#�C����m�i�+s�6����В�Qo���k�-m��P����X��J�K
�����߈w�Rhn�A�G�~s��$��y��`������}-�ǩiW�7l^���'}�O����p��ix�f^`�VM�ÛX�J6���2��B�BW~�9�G,����j	��/M��������kM}���Ց�U��'�}|���]D�)�����y��o7�~C�4ٲ�\W���y6���V�_����$
�����Zy�����{��q����� A�m�|@\�q�;�P�4�q��$׋��E��|!�e��{ ���
�)(�0h����*qS\URs�`�	�SG��?./�(�f�W��SR!��H���#�n��+������b��:�JV���v�"������2�0=E��T~�%E����l��N�H�T�T����?�y��ks°�蜻��\����P�|��\����GZ��P�)�6�>�/�����΂#�R��3�E��&�T�վ�dvmP(�#Q�)��s��c����������o�~���2�L[Qd��'��[���0�ah.1�ՙ5�!�����P�5��������jǡ��fW�yB������5'8�.2��`6զ��G���2����/�>��2P(�B+�jy�n�U'�v@�/�Zψ��S��,�+F�� ֖�6��S2Aoj���j���(��`���ICQH6}9�'t�><�2�B�xp�xh�zѐ��qpk��*�Ĕ]RAp�����=�Y��X&%0��{g��
��G��^���O���p��{ݕ�
�Z܄ ٸ����w(<odii���"��?��`��G㑅g�ǭ���:8�s��]b���M��b�l��,:�`��)��8^�p�ef"QȞȘ�|/#\��GNm�T"0}.�q�VA]
y���we����m���g�:���j�v�[��t��F_�k���b�[7z+	[����Dv"UH��-�^O1 ��,w��"��U����,}�uGp �Q�e��r��R�����H��
_���+5��B�	��������h��j]��?��-�	���m�C�W���z���� Ơ�ݎ	��b/��6�'Ө۱��&�>gŮ��U� ��<�g�R�t��yU����_F����� �,�9�k���zB�OD���- �|��D)$���Bm�yаBK��W4jj�j��C���c3&����)�t���~D��xeʬu8wv:�*�9��\��Y���X��5�%a\��*q��
�����@Z�R��0te���|�OX����Z��Y��fxX?��|����}A�`�Z��~�e7Σ�u7���`��9TQ�����m�=��mɾB�J>�lo�?��{��;Շ�W�
������!�??���Y�9؝4ﭢ��ԗ���iXmk���t�
����7wZ��]6���'W��LةK ��h	��A��x�q$�2)���"�5z%#Rf�Wh��a�-3Ɯ�dL�V:JA��&�FC�b��|���l1.�ɍꯚ�wR��&�g�T��{�5�z*ޞZ*ώ�
js(�j˸f�����mD�GJ9>�:<;����pəI1W�\" 3�Z�q���q�#q~��չ*A�"�/�h�@�/л{x��q�v���dN��*�sJ��3@w=�ݰy(�O���B}��׷�Ƀ �,q"�ZK���ޛ(�����j"jI/L��5˓����|�:<����񞽀}�#��O����A�|Q8W[P�H0U}����B�������[x�e9�&4*� ;�9������{Q��ޗ�W�M���ɕ ��M4�`��j���?Xs�/o\U:�R�5Q�t�<�d��E�+�+���~�����t��W�TZ�>.'�x���}�&P.����k+�$�i��3
�|I7������p�ٺ��(3q���y o-������� V8�0�E��vi�����R�ߕV�s� ���x����`�'��R"����5`��ʷzo*)`���?��C;�l�V��<̤WD���O�2����~�(�੄&����<O(� �p��k�^,C�R<4�����%-'�,=�u/�k�猂:�}֐�a��58#&����a����=Y��S���;�
�w,�+t��ڊ�K����B��r]�>�(�����M�ޜ��U)��?Z ��%,�1~;G�`���X���1����$~Q��53�WgV�넟�3*2���w�*t���Hժ�Bm�g�jv��N� 7�S0t!�>���i��Oڛ6%�� W�i�b��!v�	���k�:;k��G��~6��"��_ǰt18�~��q�`�����"�׭{�����!<�~ްU�`�u���P�zn\��p�Eƀ1�\��y�]þ����n�,�!����[�=-��D��D'�p��2xT�gČ{NX��M�Ջj��1��v8ڹE��IL�z*�V�Vs\i$lR+���q�F�;���X|����D���:v�N1����%Ok:��z`����96X��\�����4��/09���>�)�>�(+'��K�ſ\����v�S>w*ѓS�V|�0����\�k&O�-������$�DY۲Xa4fG�-���T-V�(.��g��,�Zy�����lh(c�^�Ӽ��m�{�H<}���3,��mIp�S�G��|d���E+���wo8KWLF��,�j��j�;4[@��_Z=�N�u~V�<u����v�R��"8z�F?fD" �nE�b�j�>f���-@rt�����X�U(�i[ɦ=���gZ���C-o=�Ag��i�ԝ�d�����ȧ��y+Յ��f`�+s�WeQ��X�$ˌ�8����A�h�9�ĳ�ָ��=���'�󀊔г�ZB�y_q�Z@b�1Iu?�����4�S�C!�zg�@(S �ސ1��Xpn���K��9�ϛZ�U��M��G�f�5z�DP�PX�1P��o�M��<A�%\'Hb/��s��*�� Ta��nF�Ej���8	丰p�~�*��g�����|�B���6H�>�����f!���'xV��+/�̟�o���B#��r�b�w�8gEA�ͨ�Z����F����	�a <�w���D"��&c�I_O(���+w2��w��=CQ�Ɛ]�"�fʮ�r�@��JC��l���Kk�x�K��f������FeP@iL�!�)q:tFN�Kح,���|�/���5�F���<�J�>�]��%��OS���	�=���X��n�ozxU�w�̖����o/�·- LԄd�/��ӽ�-�0��W�k��ʞ�5@_��B�/��t�&���,o�ovKwy"��5�<��X�r�px�3�ڦ�*���ݜyCzq�儬��d_z����!�&���%j�� ��rԁ�]���!���d��7���;��.�`��x�k�p���$
��v�\�?Z����^/��b�1������m��WEk0���.r��=h0 ���_M���{�.��_