XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��d1~��ވkT�}��S7��}|e�9y�89���B ��4�5E�!}L�OB�ԕ��<�X��gyMb�p�Z��͢�~ۊ0J���۳�uA8�ښ�ǟ�ƽ��Up�� )��}��"�γ����ޯ�Ly\#�n�\�@����Q���!��X�E=)� �[u�MIiH�ɂ���U����ka�{��1{�l��C 	���>w�s��Q�Q�]����|�1&*c��C��!���c4A�锵����z��l��V��l7�S��V�NX`��[�S���Ld����B^:�t��N�K�H?� �Xz�sa�@k�8�#_F[�He����"�3��գ��wh�
�s��y��ʲ_ j(���>`�*��k�����w��T7�(�x���h��m^��&=D߶�'*}�>�/�Eho���Z�D|F��GⅩ(�{+`~��b�T���n�t�6���_t���5AĒ�o�rB�ܼ����X���&b���,ƈL�aO��`�ڎ��]E-,9���v�tX��r*���|�B{/p3���jZv�����H�g���c�a����Z��')Mj����"���n�`��F'�YfU�1�[vJ��3��&]q
��F��T�;.9H��C)��h�u	��Ƴ%�(�B�мfi�����m�Ul���L�����
�.b`���-i0�'����X��@�:R�s,�ݢ(�Vv	N�_GDyJ���I���c�=���.%��|��r�7��������D�Į�XlxVHYEB    7744    1780I� ��&y33@륚�c��S!��tL\������Q��ٶ��?��w�w��yv��Ҋ,�|�N��߼g��#e �@i�*P�SQ|})́�ZI�硫�=����	4gH�ʯ�\9C�{��~7��Z�J�,�T�U�����]�\E���}2Qu#B�C_2X� �z`l���^�����y�P$j"]j�O�����73̣��}����I�͒H�p�9��NL��Í�:��:FC���>BY�Ogg��/B��?� c�,���ϔ��P[@���x:.E��V6�dJo2;��ǯ��Fp���d�����)\�&�-{f�:����4�%���᪸�������`I����b�!O�rk��QzdQB
�< ����֛��,���	�=�C��ln,pT1*�P��F�]��D����,�;È�#T�V���S0����ǟ�{��C�c��k�3�W����jq��jQK_~ɉz��u�)�L���[�y��V.,=�WˉrJ��3�	�<�K͡�#љݿ�����x��v��p|�U*���-UP�_a�OzP�H{�������
�M�<4P
��Z����9]��IŜ���n�%�yۑ���VT8�<!d�!fT�.}C�o��wmQ�;��x�[�'����Y���fY��V��2�0OZFz� <��?��h>��>3
9o�%����-����b�u�R�;M�.*tC�e'�|`�Qہk��ߺ�2�E.���
 '��W�x�n�v9�m��y�d��Db��${P��PRW&}��)^��+�+T�f@�;��i��$�3���kρ�Ͷ��b�`�$�F����Z�n�t�1��g�=�s�3���6�#��ڨ��g-�mȯ`�Hy�i���gT�voƜ4$�Ɍ�-���aM�8[{&�D���,���v �G���Uo���}DM�Q��p��w���c���ۤ/༰gk*{f�vG�G��P.
sx`�����{�ν������t��׉9��"U1���J�:�"��y+�q�(��ʣ�sv��2��b�OQ�d���a�\
�r�|��c���aژd����3O��ψ�W�����YFðm���g����߁x��1<BI%n=�o�c֤f�I����0{^�5��\�ɰ����M�$��͈/�,ju���VO�sFo�"Ex�&�F<�H:۟3�/A�k�a"^��Z�2�A�o�ړ=�S�ZL[����m�PuwB�6�Cd���g�q�Z�4?U`�K���Z�A1��K)�����o`}�ʶ�6���+[���M!��k�{�4Ԍeb��zi��V_b9���i��V�)�l��T_ ����"��0�3��"�d�~b|sX�TI�C7>G=Y+,���V��$���Hu�nr�wP ���шu/%�;�N��`�J�?�8xU�P�2%{>�ق��9~��A��JD���ߗ���WlR���������f��b����t�מk����ԕ<�-��W��B/ڝ�{xC5%�Qn.�n�Ȓ]~��\(dTY�stP�:��!	t������`S�G���Y���A���A(�����pQ��ْu }�Y�|D!���Qdw�f�(�59��35U7��:BV�cb�~�j�1,�d��LhW$䔎m�<~��+��;&"����D��iTӳ��R�,&�?�>�u�X0;drP�Eӷ�i��{7�/�ވ��e�"~�PI�SMos
��������(͍�H&Q�C~�*�fx�T�h�s!��!:i1��t�J�/�����Ą���>q��[D��S��W�5��ب+II�L��aY^�6�+f��"�(��c�f�b�̥��f�gzt��x�Dp�!bњ�
5@��gO?�+g��Cc!��3��E�+�=_�*Q�^ƆrE/PǫQ�`��W�S9� /�߄Ά_�9�N�M���"H$��+��ݐ7G�qB���Cʿ�֙%?�q�Ӟ�x�r�l�z{m*�ՆE�#j-�>�JASK�G��;x��ԃ�Gtd����WpҘ�p�L��@���^��YoZ+���≚�`$�`Ӧ��Zø8Q$��$�Oh!a�:�e�5�:1��� � r��ʄ��T�͜z��p��6P��(��p<Y���қN����"&�ox[qz��nءi�G�(-��*v�rcd	".�<����":�^�\��U�gH���U����/ϕ��@!�S�����i�PZƭs"����#�݁^־W���E9�� M$[%y��8G?�&�&j�I!��a��v,���	�� ����, ���$�U�����r���s:���}KW�����Eo��oH�8�#>2�]�$%I<lfj�Rp��pG]���-����P�uL�Q�T���Fk�i�`�j�a�X�s��1�j+�%ɴ��w�E�K�w�8��ם��PF|߂s�G��	��e�o�B0s3�(�~�^0�I���.�C+��[�16R7������Y�x���Y�8����)ν�PJ���x��ߕ�M��>�,��l�(�(/�\��606�=ԷC'U���"E7��Q�0qnͽʝ-[;*� �v�D�NF���������lP��4�»�W(���$>X	W�=|�8;V�c�/���M��=���)���pMõ�~���gl�R>�Vo����ū��t��7	e���� �y6�s�,��1=g"`qRX6�����4*����=��~t�R��v���(��z��@���_ۥ.X���iw����y]��`�j�"�c�W�A|��Zf�?3�wtu{g�"��`�?�#�}�:�5fLL��G�re�4����<�f�"�k+�V�����-���1+z9�,����3)q�r�Q�����'��ΥH
�{�UD}�1 Ē���p�;=�b�>:�PT�%�9���c��?�6�	�r:���&��۲�\��t���a��j�K�� R�3���0�1�P<��9��o�X�,b,�E��L��y;�6/b�#%I뤼>U����?�n�9=cDi���� VOmO[".D����g���7R���j��r:�ǫ6{�;�:�q����� m���#7����"s�W�y�����:�m'?1U}sr�I�v�%�x�KpE~]�'縍y4�u kE]G�����%^�<���ע��ėX���, -�(����m�\�ߡǐ�C�c�S�B���/T~�����ht����W��ް�M��_�[g����,��6'��PR�?�w=�ෲڠ�N95�+ �GΛ��N������NK5�icU);=�e�7�Xڲ�=|3�������x+�g�<H�i�Ml4��1�&3c34d��IE��������ϸ���~��(�=����O}D 2���K,l�%?>a��-��vRp>��n$�����&ب��N�Q*��u��.$zl�Q) �«���qލJ�������I| !2�Q/�$�Ԏ+<��ui���q�}�Da\����^3�G�hׯ�]G��S���ǿ����-!`X�� ]!Ow`��Y��<���?��5-ov>�C�����.@���eg�w䗴
�TaSy>|&֒د'(n��^E�"�p� S�Q]����쨹����-N_�g7W�������$���C��?���g[�M����qa~�+���FҤ�GM\?F�m�.�i;�*���l���7݇�/5T^q[���7�d���x�:�í���5�Bs45&T��JY�7;s}�^�H��p��KC����R
���h)�?龞�[��[�}@z��5�~��'��5�؏qՍ�[��)�H쮇��V��a	O���7�hM縳<Ɍ_��c0}���@� �_�6\[��0#k���5J�C9���F�6�K�]/���=�zO�]"�`bY>ܤr��ac�Q.g���h�2/��-�B���M��J�|c��V@�i�����3�_�@&���s��}�>85�s���2�|���\����A�)�ӟ��.Ó�1"�'�29}��,���B�T?a|yzn�ʽO��
��f��lkyt�ê���4���>�6��ʈ>�$w�@Tǜ�b)�r��4ӝ<�{�f8���BA�0��@ΈS��J3ǧVKK毧K}�l[�)���0!�ns��!+���J�ÛM��$��VU[�܏����1����Ⱦ���[�:��y����!|�X��X�\�c�^�ȓX&<�E������ޜ�)�֭�޺W��k��9v�g�2Lz��:"V+����z�HC��a����<������7,2=o��v<�$�<u~^�����Ɇ�Uҝ�T~_<�d��n(��Uf]I/λ͑I�j�'MrKx7�3�4��� �M�Y �
����;q1�6�Y���(0�]�eۗ��^��.�o�|=� ݯ����_g�`;�,u�v��N}�M{�nFHڇl;:Q{���ܼk��	9�/�~��۵��_��r?Ȃ�٤O�Ԙ3���_��8Զ��r����[�|��KY��%|�V��#����0�5E��Y�g������%_�٢L	����#�� �$��X8A{�<��.��C#H���L%�#-���� Ⱍ[���+|�ba{�'9�5�n\iEU�G�74˕�s�O��&׫@<i+~p����Q.��U��<���F�J)r�R��m�je-�)q~�ᦿ.�L!����������hp����ʤK���
�?ZW�W���`*3rsF(08G��-� ��ӥV�1.����KcY�l�1l<!�6�#&�x�E��ϙb۽��7ބdd��S�J�������%�TP��4-��_ƌ �.,}�.��O�f��*�Ɯ��va�P�i�m���N�}��n���{>N�;�0U`�=4���}��Zyt� ��]�ԬD96�n@w�}r ]�+%�����5y�������6?r�IA�(����&z�Xg��M���乀��~&�k/�,f�����-�P4���$�w����H� ŧ�I�ֲϵ�հWN��Er8����$#�����G�_u�'ֿ0K=���&3��͛�3lB�u��B!�*Pw���X��ֵt$
	-�,` �p���	X|��(��#7%�qE���dWK�#x=�����F��/� �+����ln�$��ds}@
�jA�T�Y�!-��L�?vZz���8���NA��ԲиS�y~������՘�$�!����{#�Y�c���<N�U0;�r0vӵ�z�OR��@��L8ҁ�M�?" ������.�@4<ě�p�稱oI�Ջ�jIZV��}���E܇�h�긧��&&���I�*��`��RA��D�����D�<Mo�޼[{����Q���(����^7���e�L3�8�27_��JCI�Ipp�7A�+K�O�{�� ��ޢ�T�_���>�_��`Nҽ���c���l��*�>�)��r�s�ݵf:#e�ɘta��ϡSM{�)�U��Uߋ��T�C\Vo#ƴ=� ��OC��;�fp�Ⱦ�`�z�2j�J:ϕ��]s�з�3U�$�����bJ2�	��yI�<�������-���}Cmf�{Y���?��9,<� _3عB<�#ۖE��u�����sp'˘�<H朐��ڧ��紵��Njx��S��j@�����-��ĝ����&�5^���s�S�MA�~�[�!H�c�;�CNX���Y!K�n���z��N�^B��mP[����Kc�������6���RW볿�rԹ_��uqx�Z��C�a���u��Q+�����fEc�ǵ��e>ɬdi�R�I�KxW����9Zjpˆ`ݾZ�A
F���q�h�ө�]q�e^�$f���ҬI
i�/��{���U��M���<����G����������e���