XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��W��P*j�'w��ѵ��ixGJ����:�^{�e~�6� ]n=7W�qJ�X%XV�_�%i�������J��V�Gz���"u���My�۪���� "�6>�ֿ���dOa�k@�lK3����s�ΓW����e�rA;��(��)ro�8�����[O/F�@p�Ƨ��8dcI��;qÞ�H�N^���c/��Z�)�D�3�a��}b�E��֤�o.�`�a]o��9j�����!�a�O��9��s�k7*�{��>�	�|g5wX{o�k��a��8ԥ�糍�(�x�_0Wi�e�MZE���%�N��}R3R�k�&5��m�[�x��0����&�WO���W!gT�E�c�$&9D�WiJ��r��_4?,���π�f�D�R-���Y�81��]��\G+�)׾�KL	�x��hx}�w���!݅�0<?O�,Bd(�L���8!�1[�J�xm��KE�6�6�h��L��\ޫ_j�D}��L3{����X��n�
X�?�l6#�f���BP�If�9�D/� �v��\��	�&"�8�*4��œ��g�d]��ZFg����$3��&�A��˔|8��J�O����t1�ϒ��Q
G�
!e}��o�����c���8Eq�+�[
}�ySC]�+bE��£�Qz���XU�4�oI�v�#n�7�8#�w
3���	�m�N� ����$JW6�~����)`�2���I򙢚r������)$��h�̂+�o�W���i�	�xm�����XlxVHYEB    4089     e40k<�H�bkgXU3Ut��s����\,A:?�5��	�nc��ʥh�z�_�*��9��-S&�`a�7Ҥ�5q�ǔ�/�����������}�/ R�E��P��x(@u%$*J�n�k���-��ؔX�e�IB>���ЏF���a��[�g�1�T+���� ����!l�����,���Cm�w��u ����f�����p��>:=}я4#ߧ�1��<�2E�JG/��|垕�
|"�}Ѿ�*�M��%�C�H�n��S�Vpt��~�n������E����HWY�K��g�_���
����z���j#�����e�5/�6�x�:^3��K���K:V
��D���7���(d"H�3xy@ �\��q7[�%�TN{e��0���o�h>P��ӕ���Z�v���j�g~�2h�gg��@��H;�Ǌ�p��f���[��/q��h��� �`��6t|F��ETG�n��쾌cr<u��M~���U�*���Hn@���5�����<��㡪:�˲bҿr���(?e��y�+M���i�@�ԥ���.lZ�?��0��g��b��AK7��
�Gۋ���2L�@���B� Nl�mJ�zӒ|9��+�}S3�ܘ�z���i@�w8��ck#%���8<]�����U��y��J�\ˑ�ѝX�Qΰ�{Sl~� �q ���2H�g��ˮ�rz6��"�c3��%czx�M�DiR?N�B�.��1X ^�?��$(�m�O2��������';��/9&r>xP��z���õ��s#�w�DW0�4Y�SV���`������:O4k�U/j��{�����9&����if��MtD"ꎐԱѭ&�e��_���[�����0A��n?���
�֥��^R	J�V>�ڊɌ��Cj �/q䙬��BR��8�1�X~��+J��P�R�p$�F_TՐ��D��ۆ�ϿT�T�y�k�S�L'*5����ɜ���u�E��+K]�Pġ��M'��3�|�Z�a:��N�?6�QQ��k��<����!W�vi���Ǻ��-c}<�g�bkH�-kq	�>���7e U�C<��0�(�ж<�xN>?B����79]�WaښoɋЎ�(0Jm�`�"�-�%��8\�D1"l&�s�-�����73G&�������Vvs\�[���H��́���!}��:��UQ=�!g�<�n�8�j��C�R�����R��w�7��>H$sHb]ۻ�\3���;\��O>.8i����h�U�b�n�T y}��sb������Ⱦ]�X�m9q��W��l��%7��l\.?�=�m%�w�����H�F�\��U$=#N%,h�f�!��P�un̺eP�W�4��SU�y����X8�h��X)�{5/<�d�����Zb��=~Rp�;	RGWM�v���o~C7������zB�!�d�O�~SW��n��'���OOw����K�?@���*��M
2�Q��������!P`I�z%z����9=o2p�W�:�bm��,w`a��o%c�
��lI�g����Y�IDP-ʑLW�)�@&���^?�>_�S���]�,�+m��h�֓�#����l�ۛ,�M�(���㌪�������*CƋV�"�Ws4#PXd�&�h�@
`�(NUǻ�s��{�As
�.^
�[�cS���%$G�H��i���P�3��u���㸙v���m�c�����OQ���Vq����6܍��@��"�`�x/9w�-�Y�¸I�Bx�S���H��]V('��;)Lf̌�^����>�����k���G��
hv3��n?='��njA���*����؟|%�m^^n�Є.*B�����[x
=�)B0dw��TBt���<Jw�RZ،U9}�-;:�#��gL��ߑ͌ӑv��Ȕɭ�` �;��ǂZ�K
�ؐk�����������ٗ�L�|`��誨l�Ռng��s��h!�C�(��JM��f���p��,^)�R��I�Rµ]��! ��R$Ff�y�?,����dv�+�I�W���'4R
��06t��FX�~=��*k�HVw(P��w��Wi8~m�@A�=�XLռҝ'���,��Ĩ��TQ
<��mN�'|7wU=��I����N�y�������jl��@�>J�NDt����YP'�~�x���I	��m��{����Ʋ��ۧI��0
�)P�T�S#?ԜK4|#_�X�h�OR�d��m�,��S�ٛ�gm ��>�/;�ay�/���uJ�!��k
[1�ﴄ�A���օE��; [�o�
ϧ!<�{�D�?��|G��fM������r�(���U�%܎}D��j[���lQY�D9K�:{�����G"z��U�BƐ`<!�燹��X��5��a�5��v-wj���"��*B�M���*^,f��KK8R��D�*�������ϻ���mT��L�B��2*SV�1��Et�,���\W���F�	H��EuLW������8
����(����;�\��(�"3ْ�]�(���}ƹ�D#D-��@�+��W��U���U��B��z�'�gCN����/Q"[6F�.#��x�Xpן��C��}]=��q[���a�L�H@����<�0H��F�@8Wq�(
�-�nM��Je#��x�Jp� �'ڡ����e�z�*@���ʇY_�A����W�q!�xqX0�\I���)%/׏���C��d��h�����VUl��Wئ3���%ئ�H��"��5q��1Hh��t�b̌ �y�dP/?F4S��1?��Ɠ����0\���m�{��\�[�7~41�t�syb�`Ekʡ�L.�lB�}&+��l^Ө��z�.�p<��3���ѢLi�+�F��^���^�gb��U_ZUD��/�ђ:�� ˞�{���+I�c'�V���S�f"t����2x�x���� ��D�sz�>�>`��W�A��u3s��'�5Q�s���>�ݚ���D_]^�})��M��-�x�o�b"I�r�y�Ĳ\L���X2�=3�T�\,�nÜ���0��/�΅Q���Gf��&4��Q{��~f�.{��i�x�x�!\�Av��[�R��8t�o"��5qH`U/��m�O�W)�yЗ&>�V-��c�= ��C �ƽei�2�*�L�ת��6ceF�6��� _�w�.�DDl4T&���|� �?�RZ�SS+󩙻�\���Y��Hct
&I���cRU����y���_��Gd���!��x���T�� �}��������FwG�ߓ��ƪx���z̸�J7���p9���z��^��F2����(�8cA`'��0�ZC�����{��Q�L<Y��묯>�q[����!-��/��`vmV�w��̬&��8qk_k�F�a��o��T�)���A�${᝵�<Q-�Fs�׾.��F��tV�jU���0���̦ Rÿc�[<�d���9��A����t27@c_G�M�L��큯��{��p&n�a"�T���g�Hu��%�CN��k������O9dj�w�?� ��`�S�D`�v�>w��RZ�epj\�\~��u�t�~l��m��)��ך�z��-��C����4���9S2