XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���G��$r��V*����R�J�����lu˂ze����L�K �ɞ��:�x��7�;�T���;�.,+��L���0�7�%K����[�~�Q͇����v�vo��ݬ+w�|�u��/�����5�l1.�+ �7e��y2IŤ'V��pT;'V�{A���4;cV�>D��VA4q �������)�ni}ڇϯ#��Q'|�e� ���+�L�,Xe���!�LBF	��D��1
rϐW��m������CPm�7���K+;ɍ���
�w~��
��0��k��O>~�V�7�~˘�X�G�*�XĐ� ���N��-�w	L�\�m'+��4���k�12t���P��@��Wnp��U��m�y&z<[�x���">l�G�	��'�)i����,D��+w{�Bͽ�S�%mι2ח�2��j�ޝ��ˤ�����R��<F�+���[��svd�}���'F�\��s�������/�AH�h�����W`.���/O,_�-fY�ў5}fW��e���q��T>���݂��L�(��+��~�B�h�A2�-8�ů����d ]�)��A�$|wj�ǹ<�����.U>��O2�(�������*ѯ�]:����F�k?w�>����5�{L����1���mf��+�#�)X^8�S4V�6��Z����ݻ�4��K,����7�·cIGC�]��O��iYQ�����	!�$�5%3���A'��syeq`<�D\�x�1d�؛j�Zn�����XlxVHYEB    2e55     b004�7�S�ѭ<�L��]xh �Q�;�UX����M	�k�F���k0?�r�g�!-;���H��X�g�����)�0������_Y7�3�L��_�2f! ��&اW0B�90p���	5U��ݸ�/���@f���͑��D�,�o�O��L�|����0D&d6��/�S���D���ڢ���&��kI���߲_Q��9���s��_��7TE��m�ă��J��:ā�^����6-�p�.���jX�VT�����������C�Y�Q��!h�I�O�8%H~�E����PKLφV�ҴE����!�D��D��/��r��7�&2���i���H�l:p��Ηnw��j��ܭzgF���E���js� �����^y�5Q���F: Ovy�l��"�3fƻꋜhO�Hv�^ށ�7Í�y�k^��7T�����W-�S��7���h?�M侶�(��8�g�䃢=��؝;���ۅc^x���P�h�'�p�����7�M-�T����*�7�Y�,�f�j�Rs�`��1���Euv@m��T�@A���k��G���b��5����iC)�����wU_sQ8��q؀d[�hą;�"NM4�$�!��a��Z�~�w=��Q����k{�*9Lڑ��7I��:}jXdm�kkz�z?�%���$m�e�|�;������6��j��S�9w+�A�ϰ�I�E��@�eC�Ԉ\'�0rR؋D9�$�%$p��J��k����q��2@K ׽������(���eu��Lfʏ��DA��n�5''V���N�� �T>��ܢ.(�m�]�3��
����m�:�𱺳�-�碛����j�v�u���6I�RK��_���_���fn�����w�Z9*C���,�1���4��!���2s[�p&��B���Ю��_�Ԭ��/�������8���t`�`��Rd�������U�������*�o�On�RQҳc_fn��h��Ŕ�����P�!��_���ph��
���d	�`�8�:�f������5�k26�N�xv�@�`k�d���-�H=�������π%u��n�Ҥ��G|���Hǫ\�Qﺻ�SR�����A����1-3XxЁ�e:	����g�6.�Q�W�<����Z��4�&���`�!N��� !2��Qw�] ����v�
ߒ-<���E��>�U�h�J�Z�c�{��;f�v!��M�������d���{.�'� -@�5���%���]Mz������%/�8<v��Z�)2`I<!�f0�'+q����� +i��tnb���yݕ�,"�Ag� �C+�m����^],c�Ǯ�,��^����
�⮛�5��.�~`g�c*{J
�S N���@
��k�2�HW�迹��'O��swi�IU��d�W5���K��	�:��mP��:�a������.S'�Ǵ�2"vN�:gh�l��HND��,��4ٝ��ow7=�#�#[����e�Y�C�DP!0���$N
H����'uo��4˴%]�9�_�vxM!>z�� �~�$"X�h܎�Ըs�#��/@&JC���U�z@0'nmz$�RgFG̋��8�]��ܗ�T#cQ���z��݌�{o�QF��A�_����Ϫ�ΐ��tȦv��|ąl�����~Ϛh��^���P��ޔ�%'UIҨ,7
�Z$�迻W��������/	� �e���l8�3�/����I5����h��BIr�eX[��_�t����J��OXY֌H&1��@��������9�p����yd���*�=:�a��{�H	>�J�l�9|X/w�	�{�`¸Ԉ����9�.�����S�}����(���I���7�k�8�4~��ʧT�ü�s�<HC�%�|! x	�>i�9��X5i2��kG�+nQ��^��+d@�N����,Xm,Aa�`�w��*cV���b:`��n>��@�9*J�D��h����r�o�W)b�Ǎ�={`#`Lq��~��Ʌ4��Ff�RT��/3l�g�X�t���F!�����}0�NOzM�����#ի��G&��c�ƨ璴_��I=Кjl����e0�2�U�vc5�6���}<���=��MƬ�}��Zr�كM���3�����m��F��qQ���
=��m"����
�� �{̰�zpOH�[O\Uw�2�##����;D�JI�����=������9ΨJ�)��2�MB����VK��p�*���+*i`k�Kmd����c��Y B��]��o01�{',��jt}�X� �����gI�'�J���/X,�U�
fvip�q����H2*�ds>��5��&���~�:&�P�2����=����LV�n�#}����z����t����e{��jd�ϧ�r�Ӧ��V��^i�B�Ø;�pk�<��홑�����bA_��N��E;�R/{�ν.)�������=�9ذ�!.9i: lڠ94����Ł���w�����MM��C�򫳻�Cxp'��"*I�����g�gK�(5V�ŗ�J���}ab� e���2�K��}Z+�- X؀ɯ��|��T	M�IonV��²õjuL�2�R4�X��q���RP�K�����x��w�ٖU D�����`�]�]LF}v�%�'b��s� H�Rg�$���S��xa"b�a�8@�	��*ά�S��Ԣ��Co)롡3�B��q��m+��eTG�~��d����l�����A����Kg`��F[6�