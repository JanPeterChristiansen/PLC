XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����T��178�[ي:欻�����VI�&�P\�v��᜙eӛ�,yQJ��;>�t^ 2�׊�/-�A�<�A��`-��&�=��"�s!@>1ȫ������n��H]�ѵ�zd�p!ǟT�>8��|�c����1��c|�}��6������6�Ev������$h�ސF<:��,g1%�©-��,H���k�T[0eɭ��Q�1�|h�Q��!�Y�[�dJ&�x=�a[�"'P��]������}ڻuӾ��WP0�s��X�*�U�:6��;o0d@���c\�����`���%{�2_\��p�q���++D)��[�o�E�.^���S�':�w(<ѽ�%�i�(Xc���'���6�����+�f�H��S�"G��Y�p@�I�wH�l�:�\�{�.sb�\�a��O��O$��	��a��4m��e~�'2����'��r9BKL�1^���@���<�
��q�Gr��3�h�o��S��� �-�Y(��:�U�ӕ���l���߫���꧐q؁m���S�5��Z���~�d\�����@j�{y��U�x�)l+`�anf'v)~f<׫.��������n�#Һ�s���"4�T�����>m�FSM�R? ň�w�z����F�Xp��s�4x%.B�/�Y�Y�5���O@����~	:T^+�CL_L�Ul	��]׶RG������ H41�ؑs,J˻L���"�~;��eץ"��7��
ԣ-9��ƉXlxVHYEB    fa00    2950�sO�AC�w��M�l��3�<;�r8�Iǥ8�V����Ȝ=,z�.�B_��֕5�i�T!�6{�2U]�箼H{�H��H�~YE�FB�h���?����v1�͟��Ns�3��)�,V�\�Vd�ׇfRCe���J<t~�\)少`���׷���$\Fh3�]>#O�������_*�_ c"��I�_�ej�^u	�7a���MC�?�)�I˪���㨡=�pipKDO���3�8d[?���V�3��w!~�vKLm���2���1q�NyE8*���Kv��~Ԫ�#t��gTDpU�[GH�7C�Trg��s'�Yl�>�O�6i�R"n�����I��DHm�wr
	�?1��(LڟD��.�nQ�V�^�:�����--�����^0p����r���N��3m�!J�v�ЦeY��N����f�/��I�ͻܨ3Md��N�s�zlQ��QUXsTVY���k�B$E&��6\^'&:����~�[߂8��Pm�� �����9l��=�P��O/RXx�����2ua�M��x��ĸu�rd�\�;��ZJLA0w�e6��J�Xu�F*��CE2���]åϝBK���H9�V��=S�Y䩉�Q7���n4�
Ϧ�C�����{XϥS��
6�2�sY���	�^���Znj��j�
�����ґ�-����n�6��@����o#�'�q�H0f�@�U��{&��{	��MM%Zl����wp�>������l�|�-�t&�X,d�#�2X��?v|���2���hYDi�C���E��PX��T����=;Ӡ�`�!����˜V7��~P/�.�Ƶθ-��F���)zZt!Ϝ:$ۚ"�c�5?��a���S6�9���b��e۸�>�(��Y_la(�L>-�y�\���(�-Lj!�?ֶeԲ��$�Xj�t(�f��*,�1w�N������針�"޹�M6ݷgZ����2P�5Z��-5�<�q9J%i6W�>����P9�%>��VR=��Ȳ"�%�[u��'G^����!�z/�U��A�	����L���o@�վ��'��k*�@�$4��
êU�-�-��;:�T�/N%�H�)�ag�r?�Y�3�B� �M����q?�����K:e����E�$�(�2��>�p��<� �hD�<��nj�qf��`�5$�ާ�D/&�:���3�G���Kٛr�j@B�	��>s�<~8=�xdhIfN"�G�\*���칟��S�lq��\�p�KYw��`��s�y���*�Y�(��3�B0,�-��y� �X[�d�N�]$�����(��,,B��E����֮q��~bE���\}��V���C��à첚��Kx}�~�/O��k�I7f�,rĵ���U��xM��6��[^��6���a���Ш�sGL>�=(�o�O�¾�&SY���8��\>ڪۭ��pN�
h<�<P<�Au�UzU?�$��F^�`4��{(6@�NK��|#
~�E�xU�Hnx��@�~��&�ئkj�V��>�b}o-�h���,E��ү5���%P�����W�{b���������xsi=a�5�FW�����?76��1��24}��r����+}�6��|�ᱞՏ�̓z�J���9���O�ֈ���T�d���$������ڊ�-W�?i��;DQ�8Yu!�����q%��i":��צ��eN���x��ՂK����7�/�娃���fX��#Tte;:����	6���qї�ڱG�C�}ct}O�����sB�����	�ƁOٯ]�?��ڬ� rR^�[�u2C-��x���0��Q�d��u��'JV��#�d(h[Vd��9����H�IT?��:����cd3�p���X�	C�I�ԩ{8�Y<a���O�|]����Y�nkf:�r�XZP��?�<�x����5k7;<t2�9;,�P�B�T��#���
xY��RF���:�{l���''N+��{"�����p�s��=y2>i0��m&�� *������Q�A�t#�v�+2A̋͒� 'Վ�I�Eg���LGDQ�7�u���@9����c����Yd�=�@B�Tq0�\��J�֓���x���~�e��H�3�׍\�� �����c�*7N�"�Ŵ�Ò��wP�4���C}G������=2C{���+!��L�����FE�����(%�k��=��3�݁�b���8��X����S����v����%Eraޝ�<�.����70�=%����osR��vD�ۭ+,�����e�����Q��P�����8��<Ȯ�9�N�8�`��������P�?ۛT�r�a���*�#Q�yq�xP���$��¾dw�q����k����d�!��=A�E��1j�Ɖ��>��®Kl5Y�,���S��8	�,�m틱n�GV��o��P�W�U-�+��פ�hW&\o��L*��@=j��?y��i���冦ى�D�,)`
9�gӵd.Us�Q�MG�8q��h���?�"IR���*��֟Ed�B�L�R�kW�4�\��x`�����$�&x�8���-�S�n�:N����ד܉�����Ο8�u�w	}l,꡴��{�����YV�E��X���9߶֑��"��j��#�{Ȝ/"?������dM.AFS�ݩ���-u�g@���_��P��HH!u�)��˕oWE��uB,�V�8��t�y��dAoU�m�'5�3j��Sw7lKm)�d^�\~���u��p�n����3B"�qj�9�̚�������1�(�N%:.�k �?vDL�\+�?�q�7-�za��7�띮��~$!��9ի����c�IA�!G���צu��hK����i	(j������h��U_/�-)y`?��D�j��0�_(�h=䑒0I�[��p2��M��$��s	�F�;�Ƿ��p@�5��@��e�W�J��ך�H6�jO}mOsvGi�yJ�#D��[='E>X�*?�>���m��,P?]Vi�����0�E"�I2Fs6P��e�6d�[���s@<���w.jͺ����8!�#O�N�(ʑU��A����j����ܟq@q��E~"���n�X���D��i�Ț���a��O���C���&u����6���Q���`{�8�P�l$>�n|�썢v��-�c�;�(�/E+���1�0�����zx�P��6햊����\V�[A�"r��qh�U	�%����bx�����
Pf�ʣ��C�$�G�A�<��i^��O�\CB9���pY��<�g�����"�Y�@o��@ަh+6�׵v�E6�|�\Ղ������OY���|�6u!��p�llJA�Mrn5��>;�jO�>�s�+މ��������H��R�i�<ƐT��E�#B+� v��;8�C��U�ݿ������$���6�s7�!%$�Y؆�>�l�C��@}/t)�S�>3.ɫ��t�G�hLA}�Y:=���ձ�ע��8g�qUȸ�L������.`%˕	�[_�|�,�PǞ�E���H3�3]���	"C���A���?���n�Kr7��D�S��vtt�3� �}�
��ږ�.x���K�>��z&�b	���My��/L]��~�w1XF4wʬ���)������r z�Hmvsl���S���lSc�՚��{����~vV.����J��e�=���u����$�򒘻S���m�*�)�_���JIƿ��N�ɭ��@x,|�V*}�U�!'�HM+�����1��!���J������#(�p��'���:��K�[�%[�>3r��4�j���e�%�B�]�]G$DDD�#��%�?������M���o���=��:v�)N�;a}oN�XM�Ɔw[8�VY�,�G��¯0�N�����V5K�s}q��¹��!5@�@n{��|�aQ�����괏{+I9v�>�*��� ׈�z��Qr������d�T���골���'��r0fj��+v�������{����~��w�䷫�4�$?-B�j����]^���f���&-q��D�1	$w�6�����F�!����/yi���
����3�8�q�9�$����wb�J��Cj�oES%A5��ȼ�wU[7��>��=C'�C��vA�(`�V�����
��2����98h�U]!�a^��U���Z��%��\�} ��wSͿ��aH�o�E���پ;�{�)� ���3Ƞ�l,��^��遻�v`A`�*�)?	,�+�42�6�̥�B$ b��ǭ#������xqP{�u�����A�����E(��{��[<��ZAʦ�V�#� :������P�-
�&��7���Hb�L_�3r�E�lFUݒ�4�mn4�=�S���ѭ4.uG+6�D�W���d������m���kܯB1Ė1%qU�b�� 
l0��m��4䢋��A,����]&�p����@�|�gX� J	�]ː(�� (/ˤ(�L �����h��4ډS��	�s�u�!�I� ɛlp��«�v���AGJ�������|�sIz*;�Pk`�k�e���G�)�����Z�f�xV<D�4F�x��͘o�k���x�q��$����47>�Zn�5������F�N�q`��k��Ħ��Õ�����USI�?k��A;�G*D,B���nځWWn������.@}��bq�(��=+����J�|q'9'��e���s�)|KI�����I�ִ�V�\�h�1��	�@�i|�,�������J�;"i�3�ڷ�Գ���&3����r��Z�[��(#k�62��1� r��{����=�H�e<�Gͻ/	`{!/AZ�ߢb���Cf�a��r�f*��P����=�S�(X)˗a:��0>�2?}*��v<@Կ19е�dP�ԉ�l���<J�\�B�6�I�r.�Z�s4�%�0�湰ٴ�����'eg�/tW���u�G����3+׋c���0��co�_�JR���[ҏ�ng�'Zh-IOo�����Y>�9�cU�����z�ȴz��S�d2��	3�pY�����Wr���������%
[�_8��~f��w�C��e���M��ic��I@�eLd��3uѯ�욟@%��Ү�,
T���^:_���9��@}3Ԝ
���A��� �8�
��sY,����#���*j�������|,��'[M缴!���_?Q��B������Ϋ3e���/�^��9�{����������\j �<�����ԃ�ף��2a���쨮	?q�<�?F&���s��w�.WM-6`>�!�jb�l�Ә���u-z췭԰���@'�����(4_J��~J����)����G�j?���\n!���k��U�5� �y.ܕTEQ:y�H�SV��L	�v �[�{��T�f[�ѽQE�a�J:Sy�絀�b��[(6�����G��W���v��������_�K�w%�sk�r�l�i��Ŷ��m�l{�F*l��/\�U��Q��
8�w�-M��C'U7�'9�4X�n8��ܦJgX[�Lb�X�:�k�*ٷ�O)r.�o�|Ӗf��B�v�/�b8-����N���L�Ag���%���M�d�uҍ���ꚲ���z���)n��~t����I^(.�0��-�юim�*�r�tYPK�[�R�X<`؉��dЦ���#'3�`n�KanS�b^<�Q�l:�L��q��H��>v@	Ϙ�f>,��s���W�w`��6����MbO4ie���Q���W~�e��Z����R�zx�f ��4��®�I^
�j5IpK��<]��_Er�D�t��I��&���cnf/���	���2��#�7�����]��D�9����l����<*e����,��*�E��r%-��ꀗ��Hѭn;a�L��9w�orf%U���G��_�5�XOv������h�T��r�D�u(>�][G���G��V�����Gp��uT�\f.q�����K��5H�Bw� q��������b ��҂A�D��C�EQ���
w[J�/����iO����#�w���v'���k�
/򇾱���D�q��ͺ_ʌP���nK-m�X<G#�mZ㵢T�pg;b~j�r C4BH�ò�q�wi����puh�i�{b<+�9jk����i�I��b��X�^�i9g��Xf	ap��s	{���WFQ�V�ݟ�-gF�8CF�B��ɭ��7�I�Ke���h*�����v��B�'��Ӆ�-�<+|��;�gk
:&*�_�)x���Ѿ���W�Lbm��a��c������dM4���<$H�A��$��]�V��_z�-׃� ��y��O?�%{����JX�$B�s*����T���Ӿ�����H�P�!���{VxV�2�U
rU�?_����g�'�c���*FY���[,�fe}0K"n��K�#���~�<�6��#\����"�/j\��;��Rq��wz�?\g��&�M$~�G#`�\ .;x?@h��Xs����:I�ۻ�2��׵�:ɹ�ԩ�E��_��%�R���IK/y'US��X�2c��$�cd����O*���m��[ܣC6��M��������ٗ)��y�w��[��ѡsQf{83IͦF���0�}�X�?z��YmΦ���3 k�z�4$�g��;,:�q��^���kHm',(�]T�B�{j��j��k�Iue&�U�<+��H죆����9#_ �G�$��J鰏�<�I���'K���:��1��ko�9J��;rX��#e�;���ѵ�����l
�R'���H�X�b7���_,+�/[\�(�G�G�����҆R��E�2��� �	�����Ϯ�7�!~��S�� f�w�����kYי�|���9����"~>�\j��O_�,�N�Q����4�K��8�N�ե�ݹt|�[x���0_��az}�45�C��"N�>�j�1�Z(X!�s�2�v�#�%:�$��X?����}�*7����9��Dfn��EM��+���7�}�"@u����z���bg7���<&Łuh� �f��L���lk�����s����Ჳ�gֱ��z�dX��=,�W�P�̧�o��L��׶��t�(�PUuz�A�fD���5����D(T�Y;4fYΑ��91�sցw����>
�4�m�0��n��G�%֘5��ؘ��?�JR~��nۡF����y��">D֋0���
@��4߈Bn�� _�A��B�Y�U�j�B��`4� vb&��w��n�fA��;��O-��9K��K�e&@&|inu��Sɹ1����я=���r�����rPf�bg����om�e����ð���U�4"�ķn�K�J����`�[�ֈw7��g�ǔ�����tiyi�x֒��x�NT{W5��$n� �EjJs��zY���ϋc�e2���� �?
t^��¶?��^@gl<�0��f��3�����d����΃kǬS�s�[�T�B+@��ik���ўD�����eE&������F>c�N��=��߹�6��҂�\D�&4nv��Ng�,�ѫ�������	�j#��v��2+uᑣ>-\-��Q^JYp��}X[.�^�mh�� ��:�������C>�W��?j�I�0���\u�Q��*m���tMoI�Iq�J��_&0������f�ډd<�|�H�g�b���F�A�ܽ0Tڞ�p�����N�nc#H��bڧ�Է,�����T�-���D:�uD�(;�d*[A���R`B����� ��Zi:�ъo���=2�4=~w���ØM�	b0짇�铍N�2*�U`s�Ӄ>�1�!kIj2�:5ɐV���R 6y�L]"��tH"���Sf�W��^;�;��R�Ú�t�P{y��5C,sJ�ˉ�Gw����b~����!q�\��]s�����*ߌ���'�h�1�'JA���{��V �"�\�8[m�3��K ?�6��N��(=4�I���a��-�Gl�&�����7r�K�=��{f���Fw�q*A�a���tj�D8�~��0n<�-}֭|xb+_��{�cM���L�|\V�ڮۇ�e
��ܯ���"�b�����Q�_���:=�T��\�%���)٭`�CIz�a:�=�I8LG�Q'�(��.��PQ�Y�U��n�0'���(�/e��^�51.���(,64d�9J'OQ��Γk��n�ڟ�*�ɻ���ɞA�G�g�	x^Bv(�(h��V�z���n9��� ����"��-z���㮊�燚S.��_��Z��'m��q\�ؘ����9W;f�'�\��$������������U�!�W�	&E������/��N��r�:�lF���n��ji�K�@t%�E#CƂ��`|�[�n}��2?��!P߃4��qLSE��I�l6)��TdY�`��Vd�@���$&h�&.��Т7˜��B��D4�R����p��*�H��f�a�X^2�"��n�xdQ�-S\C��f	��E���gFA�z�9ܿ�zE�J[���B+���e�+���M},�߯�����!�S\A�m�%�l?���0Cͨ�&�7u�SdL���Ӏ�n���8דD�{ܠH����䏾�C�*߷@ؕq��;��A���ܧ�p���B�����[�>^�=�{�ɻ��^��V�5���|�>	���7����4�
��a��3���]L�*^Z4����C<���	��洐
kw��Nz�2f��|(�<�d��Le��:lO�ߣ�e�kB�^�	��YW���;�I?l�$���Ww*�\�!�{��3�O�!b��i�$�Z�2X�����a�?�1Ģ��"jg�Pc@��N|�vE�^���� X�Uw׬?�<?��g�J���:a��~eU4��"5R:!W����ɼ�|��Ġ��J\�LI�h���cֈ�io��W�����{���
�g��(����p����@�0]���i�"tda�uzk����{�~e����=I�Y\�R�E�}�u6Wl{��]_�2[Z�t�O�]'}��f�B~®d��x���&b0�^��j�b��	���M\�GحM�j�Q0bR���,�Q�-��ظ�!���!p����\�����A��@aY?b ޹.qdZ1�Q-3��K-�
Ya*b_n=Z��/m`���T�ڠ&�ॊ���s�Ĥ�J���YP\i:�Ι���Q��%���$�Ϯs���fƄ� �F��,�.�j�x�K])C���T:�}� �#У���#O����G��|�4 �!Z�$=_Xӳ?�����kPG�91��N�����˓O������ ���h:pU.�|ӱ����=7�w�Μ�8+�;v*0H�	Xp�U��iZ0���e}����
W`K�O�m�אL���r4�|�^)���j�у`�����z7�
����L�#�������De�K.+_ݝE)�v�!��+�0�>dr��'�݁�*�m�~��ϬAOi�K�.UE-#���Q���z�T��[�\�it)������Ƒ�f��/)_�`�,�axD&@bT�kz�����9����E���BcZ��Ǣi��^v|i�Ez�}�ή�)�����O@V����B���Re��x�i�y�F�1+?&���+�%�%�����c�AxY�P�6RF^DB
�m"[T��Ê1y}Ӱ�u��@�X=H(4�#\N��`�O�c��;��Il�!h+��K+W�������4�*%6��:��+6�esqh2��v|�N���R�iVv{=�w��9���e��%�=@�|J�}�L%�1�JU�W;X�I��R�mv2�e��TWa�޳E���͑�Jp�)�7�(���h�(�Ϊ�qũݻ�\�զj�p��(t%�(aF�tkL���1߄��(D�n0�Vo[e֪x��ߔ���4?�Bެ��D�5��Z���}�1�����	&ɜ�9�M�ð�R�м`_A':$����L���u x�v2�n�I��R�%��}Ҳ�7P�����j���Q�\'�5��@�D�\Z@��1���2`/�xt��i��F̙�Ɓ��f��DHuF�J��ݯ
��(-*f�6*�;2�AB��g�1�4p�+.�ΩNQ�W]����j�	ؤ�5r��tј��r�N����!�۹-t�-q3�gP�N��J��EXW.8�������"�l�%��ǩt���Q� +O�O�o�y�a�vY�|J���s{υO�}��07޹��o��yƊ�)������Y����9�u�B�8����*�j���	��dz<Ij�}Ӂ�o�� 2i/�L7*��(�^����	�Xt����N˕(^���~1g�Q��&�=�ވ��q-R���=�mXlxVHYEB    fa00    1e30@�A����b���yN|S�����'�\b�حL���Y�;�_g;L�?uhC���F��kJn�������~��X4�P/�
��sU9�_]�:�ҟ�,�C��U��ͽ;$I���^��r�_�@Xƕ݄'c�Tp$�[!����0�Z8�j�N� ��[���J(1PP��N��vD�V	��5,���W�w�f��[ZV�������X%,�j,��L�N�	��di39W�B)3��]f05��:�Cm���C ҒMY�xU���4�3_�e0���������z��/�X�v����(���*;LA6*o];sf�z�^]6P��Gi���y�m�S�H�+~&�a�!�x��]�bI�3��*6����H�A�y�|T$�)TϜ*�A!Rv��ncʹ�����%�}��C���Z�������ҫ����x �$�L�����P�Sy6\����*�Z�Qi����#)���^/����&�Y]��,���AlqCs�tO]���&���33��q�1�MRy����\���*[�V���x�4���gJ�G4mq�f����SQ�*��!1��*����u���9O�,U8t�=I�H�^V75����Q�0��K�0����`�R��)*���`@��9��H�׮8��dK���TNp.�v�:C5.�����}����SP�R�g�����v{`�T�">}��g��l�V��Z�Z�x&��#��b	(v+�������	�n:n��9��QC2_�ڡ�85����s&YJ��͡������>g�܏xLv�t�(�=�l�ȈA��Ճ�/f���+� ,�����5���P�L���T)���-�>��z!
��HO��-�q�u?W~��C�N�N��q`��=����%8R��A�R6MN�����fY�o%Iٸ<)�K3��4���Co6��3��_�0��{So�uOCg5��� �>b�\�:���˟�ܗN���H	��C���>��f�)�.�d-O�7��ǇN�x���!"{zR�ZY С;k�7��&t oѪZ�T"3��-�\�i���O�.�^&r&k��kL:/q��r'�؇�A�p8��0E��Z[��ۛ��fW�x�ttǲm�S_��z��YQL+�����-�{�߳t��]�F$
�w�V�;M���@џ@��6�nl-Z�-Zz��~o5������<4d�4��4#�qt���t�sd��^>�Yu�`V��%�d�"ɳa��a��"�S�+��9�I�-��N���iv�y�Ȓ>x�����p�O��>5B�m�����=,����_Bg�s�1�@7\�_�ũ�`Xys����e���)ǩ8����q��\/S��N�S�Wط6�ʇ��=����f�:)�A�A�C�l�6_�@��X��?�F{�'s�%�3�e]Ϳиm��Ѹ���Y@��������j=GmKj�*����b7ո��S��
�'�����B�&3�o�1�Wt�f�U@�����i|����d�d/�*�F%�ez#a*��6�R����w62��uF	����"Z�$��F���ԝ�Z
R��6�9�|U;�#����[����Mb	�����j�ԋE�j��a�,ǺP`n=kH,�r�eZ��!���t�yQ��NQ���6,U��<���rJT�* >~��	O��l�(���)���-�Qz_���Ԋ�6��6�%����Liw�˂ⲩ�/���S�fq��x��	F�:RJ>8�eį�|�;�A{C��b�eϏoIF<����Y�7���-�3�r�~w���j���`��뽚����e�.�:��?��O�B�sL�wI��{�7�Puo����`�����koK���7w�%׋��^��}��Wl�
F3�9w*h"q�A�M�(p|�O��X�p�QLh���Uo�j�؎��xBH���~�b-$k���)�^�_�G��ʞՊ�(U*�|USU�w�!}��D�|��4�_�/��u�Qv-�ޝɕ������W�T���!<	6�3����e,u�Di�)%��'��`��Y0�/���%V�8��U���:�Z�WO@�N@�)�S	��������Vx�fs�MBOӳ3jf�)ҍ�e��J�����E�bz�ҵ�G`F������u����N$�p���Z�t[n��o�7��0��k��E2���_u�B����#�IH�/I�MT`�cӼ�e��%7���͡	,w}r������!�{NL+$�ªj��Nu�� H(C��/���.���"��D��@��uK���îQ!.b��!:�ј��{T�N�A<�vM�	��Y=PS7��X�*�EF�7� ��ޫ�Îi�A�D���7���`>�p�rC-��R(�E+�����1�;�`����BU��2v`Ua;Q�Ƞ�H���a�P8sl�_�y�b!�Rt�RX�M4Ki-�LA��N���O���o���	��r{6�uvw!�Z��A����-Pi�V���"���#j�{ń���0
Ph$�����@�e�E�}�
������X�@X��N���Q��!U��\)	@���ϰ=[Ԋ�Sc^�hݱ���n�a��$�r'�Cf�(���2g:�ܯKR۶ҕ��u���&�Cs��7k��'��i�t�_�6��������fz�H;�{�ظK��o7r����7kH��Oy�~�:�+Nٲn��otm��?Ґ�Ca(���-�H_hz����
ϝ��ɭ�L}���DCg-W��6ĥ�<���>@������"����N<�V��?� [��݆�����U�}����8o��nhB���m�[&P�B�z����ke۔(w�rğ�ٿ��W�ػ�&�w��܆t�d���.-cQ�ߕ�UQ��J�}p�v�ƛ��v��)��	1�ﺛ�,���7���}J��ۑ�=���Yg�A'�]C�d�j5�8�,Wfm}��'}R�+�ļ���D��	"�-܉��:M�u�d�U�< �}�=�L-ɹٞ ������w�ەڵk��E(Ӊ4��dXi� ��I��D��K�W�ݠ�5��a<Na�ʆ,�M����u�S�<���8%�H��Z� 3�aw��f��9|�;��!`��
�"1������W/�@�� @���e���pO��|�S��W<ϐ�8�&��B����������g4����+�ǿ!��#�K4Dk�G��}�������4����׀;s���!��|>=��27��VGǇ�<$�l]z� ֙���;,����'T����~�=3�X3N�Ⱥz�XR`!�)�r�䮻�[ɧ��os��CKD�q���%�g� (=�J�߬��.E��Ѐ���Y�����NE� ��ܺ(�pu����-i�Ϡ�K����sT��L)Q�2FmlL.٥Օq �E�7@N;����5ƒ�Uũg�oǳ6��'C�Z7nk�X|9=7A�-Ak0�x�[e	֬���r*�>z!�8xB�����-h<s�w��n�o3	Z<��U�p$�Eɏ0��k�������Z6;bǭ��l{$��\/޽����ŉD��fm�T��	v���!���MDh�_3���9�M�����ݐתj���n��A�L2���=.�B��m�~�%��
@������9aGڨn2��ve�ȅ��]áfi�q"]ʎ蝐y6G(�@Jx�bL�TR������x2���`d���<,��?N��}x���;��� @v����0��ڥYQG�Zb��Z���?��S�*�6$�M\�o��7���>�ݤ\]Q���J_�A��	K��)1�X�?k{���o��տ�_�;�j1��iZ����5{��i=9�`�w�L4��.22�ł�Ov#��q��D�H�1?i�e)�;a,�ܹ�5�T�zf��Ur��q�6B��{�n�Om�&F+���X���V�*6#U�1u�:�rh}F���vx�c$��P�+��P�Ɯ���K�n�l:�u�`J4���=#K�r�*~&ڝ�2��|����3���|���j����6ú-c����T.1{U��'&7�Ne�V�4�̱�F��]3 �ib�F��߉R�_���Џ @iٴ��=�j���ϖ�����s�=�j�������!�S�e0�C��D�s�zԖ'8~`8�L�ѥ�lH v:�j�����I��B��UAg���ѺfG1t�͎��W[���$fU��r�
v�$ C�b�Q´nQ����%Jgan'B�h��o��ns�#�V���c�
�����)� ��@�.�dN[b?4�C��L2Z3��M@|�/��6I�;�Q�7���|/���[���q(n��K�@㥋>ĥ��.��HS��%�UG�G��yKhB{��`�l��ʫ30ͯ�p#�l$B�m��Uu&�Y�VS�ǧz�:�ӛ���%��ȳH&`�6!��&ʌ�ާ|��xi��j��%2�3|=�+��#�h�k��ȕ�/��	N �g��S�K/��Ntq����I����N��S7�ł�μV0�B��s?p�ܲ�����;�nD��2�*�������L0r�����#j��q�T<�2�k��"w`�'������Jݸ�!aT̍Z���;ֶ[����.8č��BtJU�0i,�v�|�� V���Y��tD�ၦ:?�$;rZ�pb|�6�ؔ���!+�G�^�ꮃ>"�j���4�(��g:ћ����{k2��-y�y'x�6W�a˭��
�2�A7 �L:�,L��b� Wx=� ��SE�a%�&0h��}��������%�U�CB!�v��U�6OQ/^�=,�Ã��ذ���['��up�	;ŕc����u����P�`���dM�aЌ�\�\z�u��/ӝ�,N�2���`�J�',i�P^���(5�����piRS̟ и�� ���_	Y{����*�?m�h��Z@�����X���	�K}�N�3	�V]���\E�&�ɾ���0�y�8��5)��Hn��Ī��F�	�b">��J�rk�äT�۵^�:�2�\l]�>g?߹$+��ǝ2%/oK'W�&$�v�׿UVD��d53x��0����s�L�AM���P�P��L��%wkG�T��dD
�?ͭ&�N����[��0�a�$�h0�x��CQ"08���u� 9K0�nWn=�d&������q��}��V=�֌���v�������5{�n�$!�ޓWy������[�!�=s�W�
��p�r�'��[�a1]��|.��[XA����yA���HxK���Nn�_s��]Ȫ�wt��B���^c)"�����.���o�g[��C�"�C��ٽ��[g���^zoI�u �7� �Ǟrm�A�1#ղ��\`{f*�Y5�� �C7-цf?.*M��}{Y��5`' ��"��q�g�]�\k�!?��	�_'͛������2�*�j��/G�W�_h���ۄp�g�L���m~�s8ؘK��(A�2��?/�^�{�@f}�*��q��3ZC������2����X�[L	e���[����%*�~�����Aq�N���|�3������<�+�8��9��6 Mw�܉~��?Sa2�z�H�R�91XC��X�A�$�G��˗���VH��ܿ���6]���:q?�����"K$�
��aòu�#֍�L�����}��S������&�4���Rp�[���ƾ��f!쐜dѨ��T��$P� � o����I3����pD8en[dl����_�Zf3�C�����ȱv���ҭ�]�.i�(�L^Q:7����
~/�T�`M�a.�a�"@��ԍ[�y?A7W;#x:��١�&e�Io�]� 4�Y}��""2?�h�|�[Ժ6Ǩ5����<��_�JmN5�HV-���=� �\O4�Ka� ��Ɂ��tֹ����	֨`D:���}�~���7�b�����T�	� 8�G>�D� 
$�ǂ�Yu� ������t�Xk`�	��}�@ �;C����"���Eh}���'�x�QU�|߂���>�u� Y�N�r�	Cs>�;evc�*A�g�ɵ��n>j~T2�j��4�0��`~�ύ��<-����5*�L�K�=�{�C�e!E#B�%�����_t��8
�w����.�T���N�\*�-���T0�>3��A�ތ\О��<&n����Q���#����j����L"���v�U2G@��mcG,`7<�C�*���.���xv'�^�	]��@m-B��bI��$�)��{�C-.3M���W�P���n5>���h.V��_<�ǂ��f�'lB�C[ .c�o�C��O��El�7V��咯�R^��۠hu--��S�#*M|�F(���Hɳ�w+�`vB����� �%^����Kg���*��Q�	���/�eq���^qo!s]����l,��?XS.+o<��!|��Yt���;5�#D�9�p�Ί�����˅�Ԁ��	�O0��'���LX��K݈�����o\��e��6�a��S��)�s�A���������kS�qI8'iP��զ?�DS.X4���L���>=i�lT��>��Z�$�G5�O�l�WZE���U+C�#��٤���}�+,H�&���:9fLU8Jn����2����AAM��kL'�cB���n��h��M��s�'榒�A�.��%�1�L	���>� ����I"����R~�|��U�u8��s�e|!5�X�#�G/��n2��J�����0�����!����$�bW��H@�A�*� g0v�!ј�>��Lω�����x��ڃ�!&��l���:�T�,��u2�f+�AP$V�Jܓ�ۣ�z�	�������i蛃+>��6��Ө{�Fx�g��퓟����ϱ��f���!S���&c]DQ�>�l|�P��+� ���ڹ�c'�^�"�P����Ǖ4 �q�+M��8�'��,:�]�6:����׼S~���*��Z���_�&f]��iy"23C,kK͇�owk]�%�#����#��E��q���$q�J�������G��sB��E�GK��N�b6��H�s+���]��
�ɹT���xf��Ǒ�=�b���S3�DnZ�0��Yg9ն��oxt����pQ�͟�=��۰�w�$��������dZ�gg"�\%�2�5}��`l/e�@�&C���iD�X4����c��$��CmAf��_r3�=���OQF"\^��f�<�6����`IvU�h��.���C�^�Z����)�Z��]���S!R�]g��
s�����6��U�F<D�5�Q&
U��2dH>�x������)q;<BU�9���*`�l�Lqq/4��L?����!���{�pT�k��4/kƑ�}L��w����hAb�C��F%Sex��١��ϱ:����\��iv7|��K&i,�˛���^�e\�k��Y|8���"�~R'.��ؘ�����nQvH�.�ԶTy�>t�t��ܜ@�#���5I�|d�&S�sN-/�d�vn*� ��N�ףO��2l�[i��u���f/'�N�VI�VD��s�ɉ����������k�sT�iy��\�[�����P�w�&a�'a-��+y[揇O\a-v�䝿�C��ņ���XlxVHYEB    fa00    1d20,q&=4���2qM�;���_�7�c������wP��ܚ���OJ:(Ȕ$J0�,�ФF%x9|W���x�+��; ��et\8��8h�Xa��"de��8;WŞ��8Nݹ	���+65�Đ`� C�[8����m�XL��{�|et���g�����X��n�I�)L�9��ד����(jΊ���4.NFou ��ZS�����k����X`���=h��*�f5v���g�[H�l�K퓰�]q�6�LyB�1�'���@#"���#M@�p�EǓΔ��/6��W�PZ�M.��+�:��5j'�E\���2�	 r׆I�i�e<�,���߹�.�,7࣊�U8��h���=	�[�#�t�����1���Ty9�!UO�X�6*��A�ߋ	r�8����$'�N�Hز�H����(�C�_�l�ʳ_P��%�S���,P��LTh�|�	o���)�,"�N� y�5+��d����Q0�4l#�Qvm�q��ۢ֨e��z��Ctӕ���3�����pe�Pr �o-0ewu�ı؋�ζ��Z�KO����3��jw�5�T}
�N������+9>��̕r�!���YZݾ:��8su�z���-�KT�?�!�T
.+gn��N[ߨ�Sg~҅���\��b�N#�)��&-/}�����5�����s�k��_R��:�j	�sw5���u;tn�t&@�4�JFM�il���(]��!m�z> �TN0X�b�1s�H�����
�`7��R}����G��npv,Tğ2֣�+�(Ca��·�k�&��������g��h�:�9�eR�7���������t4]�A���^hX���\�0���� c��J��Qb��_n�������^���%�jc`Cn�u߾�V34`S]�0�@� �QB0�Q"�1)��m^�1�.�L�jW��)v���@zNa�:E�k�g�o��̵�[��,�5V�Ǜ�Q����rAu�0�g봰ֆ�غ�[PyF�_B ��P%%��;����vX�n�dUG��_��v +��Z���r=h��ހ�t_��6���-�| ���ۼotxG��ºs���gY���6๬��e��.T�&�4f�B�[�GFW'����K�]O��[(\���zWmW����9uM��=����T�������"�5D<[��w٭��y�VfR��ïZ
�wykk<M��+a�@���$�YX40�ݱ�d!��K���|lB}��Mjk��"��+��O�,��_s�C��������%S�}4��"G�~�kz*�W`A.�5�l�m.1	p�ŽC�vA���Qw8XO���o�����M�pS����_5��=yf>#���}t�8P�_~���(�����䘒.����d�� ���r��N*�*\g������{1�g������x�M���WI"�k?��|��]����6�!���{�'�]Q�C����V�q�l��0�l����d��i�F&���;S�kj�S�b��K�;E%m`L���??>��[��.�TkłF �s�P�=�����̊��Qʁ�|1�o]'(Z�1?��[FJ�������i�?��Jk�86�
�"9��q���tWܮ���8/�TުOS��7��l���m �+ҩtm�0�����]���<%E���a>��ijuV%�,��3�n�Q^�D^��/�4m���~� ����~��PgT趈aآ�t��8�*��U���.{�����sl+����N���;l�l���y|���΀��eu��x�nMt� �lQ
�!�@kڶ�)�[��o9�����v^���tVg������(+̽7;a��b�>�\�o` ���$��b�S�
�F�V�WT?�p�4����2����6�-C��������P2mڑ6B�����Jup붌��1fƎ���L�ZZ
&��Ġ3E>6���n��*�yX���?�3��+
��@lJ����i��o��먉ԋ_Q2�(/�z��(�#:_��>�S���^�`��Uj��Jk�]�J^�;zt�0�������u'7����v���S^����_���dnh4m{��[�W�~<f�=<�`���?�N�� %;͜��?��"�&k�C�u�h�t�/�L�q����"���H|�#-���Z�/�h����t+mr�dp�H����!�V[��	�X�J"v�!���:�J_��J�� D':��w�\8�r�Gvu�O/��GU&�8~�����X9�����I#�Ҿ�C���R}U����|W1T+��g���:>%coxu zX�j僿��W�h����F-1_�_k5"	>������Ж)�5�l�K%�����V�W]t��(f>S��N%�G����L��~!CP��4�~2^��`a�8���V�$
��Q,Rw]<t�}{��r��L4H�x}N�6}'[�Y��m0�>
�X0�ꤪ�]w��v!֑�_ii��T1ד�%g�A|����D�a�����-�VJ��k���rٖ�ƿ?��?�،�*Z�	�6N�9^~C�A� �E7�`�ӒH�y"��ax�e�a��I���K�>�I����Lo����#������S������rц�Ǖ��t�;���$�Z�v(����שx��wu4�Ӭk�c��̶z���r'jwY�0���eA�L��zpm���/s\$X�r-S9ݡ�#Nok���n͗P�HNka�`�Y��J�gk�X���@E}K���Y�;�r[p��4s(\%��J��:������ʜ�,c����05@+|1��SF���Eb��J'��q.uވl�)$j�����{��a� �)Hk���-��	�X��Y:�E?�(^E��}�B�W�;`l�Ѹe�g�O�����1у����Yp�e�ma� �	+��P
i[A���G��9-�nލ{�<y�y�JU�<Z�]d�x0䊜�����7�����?��^&��`,J�*��ϯVO�9]>�@=�����B�N5�`+�w�-5������3�|�}�qA2��;�p�8~7�����I��ϴ���o��_x�P�IM �&���W^�o�G*��WD�9��e5h}��N#�YE|���1�y��C�`R��:wG���d�Ӈ�S�GN�#�B���`u�]��2%����"����R���sZ ���w�����&C�w/e��l��q�&"��u�:	]
�.�]���;�&A��8O��ڒ �Pݳ'��tO�h�0��U����� nu��	�q�-a��F��wVW$�Y�F�އK� B��;����nt��J*;��.Q��>�ɧ�G���\�#��!�Q����$���UF���>�z��گ�t({ �.=<'�~?�k��L̒NV��M(���9�qZ��O� C����k�ߴgc����u.������W��'ی:����㝼��	wwZ΃ӈ^2���
A��T|����=�< fmX<|��;녢�ʫQ�L�bapL���
�3��Wb3F[kףW�H�J9�o��Z!!X��G��pk�Nm�j\�q����?ED/p -^�Ì�{���x�i�h^�>Z+ڇa���h�7�x��H�VF�+[�yȳ�~�˧nK���`�$��3���Sy�_����pW>�9w����*ٟ���8�2��2 ��z� ��Y<����FpvXW��d���$o�5�ޜ�;��|� ���� �e��ȳ�Y%��\��CC��\�j�Q��l�x��K��ϧ֭x׊I�C"H�&(�;��;;g����2Dy��~i�X��"����K�#Ok�Ąs�Mm3���E��+_�ܡ��� �4~�j�{O��g+yA=ռj�C��-	}�� W�Ѭr��D�M�f�{�,,\eqQ�m��j[1be��A��v+����p&vWx��V�po�aƛ��0�yC�<8C�h��4E�5������|�*Ҥ�������L�O����d�sx���u�-�����_�dL0��g�(�{��&��<�5wLI(��N����T_�h^��$'�N���<�K;c����{���p��N(UN�6o���o�S?{�,�g���>oO�	����C�Et׵���%Â�>=]G!���#K�n�;��3.�V;�o����r��3Q'�Q����!��]���;rlj^��xw;P����c�]y��\6CL@�5(�5$�����l������׶�����ȇk�xL��9k�J@ݩ������d���<G^���ݴ���. ��z4�R5܈ۆ�0��uO�é��p芓k���v����hf��4V2��l�L��Ml��ĳ0D�@�3	Ŀ��wm#�Xh�G��^J ̜�y�{��`���g~�S��F�B$���#9���wL��_�N�R]ɡ�Ơ,�ڥձ�p��e�ehz��|㝮i"�7�_�Y>�O�7X��yH���>��}R~��V�_����JFH���X���T��d�I:db��&De�oA���l"5�[�8�U������w��
o&����$�!�P#�{�����z�jdnb�&%E���rʂ{������!�3ts��dӫ��ܫ8���U9��� ù
�_yL�v�D5|��/y��f�iTh�|����P�C�z"�#>"�����e`����pc�_{�d���/A��x8�p� �-�qFծ���� �;�ٳ�����G�Rr�@^Q�c
�9�Z��+���C���l�pl��3�>��Ii�v��qa���B�d�0wĴ⫢��K�+(�l�ʪbcxip�0Բ��ձ�.*I��ZH�P@��W墶l�Ѣ�V�SvB�#�Jb,y�X�9f� �l&d��,���#�W/��]���X��4��r��Z�l��%*�Ug��|��1H�� �7T��<#�l0\�<@�[�A�V�,�H���*���NN�}X��eǗ-3 0��z��G����Z�|0�w�6�d�HV��O�<���!���`K�0p�F0�W�������<Q�:LC�^�RE�d􁳠�Q��t�I���b�4��� JO��]��'G̰�@468\����v�T�lb���B�����,<�:?2�1���#]�-=�tਡzPY�]�?�1�=�^��֣����.H.ݹ����;���t�5)�W��'��3~���B%�/�9���ٓ!}��S���ێ��)FpM�FD13X�՝�|��Y	��kC�U-��S(>�������!w~���z��g�a�����A��V�7�fa뵨����U%���=7��l�FOoP�l�_^���8��!N�n��G'J[v��K�߅�w�/�ߊxn�i���I +��|T2���<�fO�rs�gX�f Q~n�T���Pq�����O�lå�jn&�n�:Dd'����e_��S�(쁻���ј��N<жA���9G��ҁ3����ƈ���F+_`�"�_,nܷ1�-[sM��������� *|�� �j\nu�y�65��N~F�P�O��mA�5�����Ol�P���R���"!�]���A���$��<B���4/�C
ϯd�ҋ�=�5�x�!	ҥ�Y�'Q��s��28�)�i��_
��z���C�����R����̆)쀎�� ����^�`��|9�s��3�y��%����}F0C����~���j�r!�V�%�2��aЮ� b��z\����w�<$��/9���{l��A�H�����t�a�75}u�F���\gr[����*�F��ef�
|P�"�ח��Rs���x��w�DҰ���e��s�]���9L�<uٚ��CsCSP�e깏�M5��s�8q��n������vf�&��:I�d@jL������ig��7��%_�Y2�V�O>�@�a� ��(��U�(�0}�#!?}'GuΨD���j4D�Pi3��(�xX�%>rQ?��n�Af&E�)�i+Z�I:�U8̮NY�N�Nܼ��Z]�_F�Q��^�R%�����ϵ���8<i��q�1ߥ��K���}�NeZ89�%��?%ѧX���P<�
vy�vЗ���j�\�U2x���B�GQ*]�P$�K�i|���2�l�����Kx�l�
��k�~j��;p�P�F�%�����K�j�>��90-���`&��V���	�ώ;�ɌM��AvM�-�N{jz͖
Z���h�ӻ�ڽ#�1�UK�DT�wɍ��BI�B���q�n$��L,��ڥތN�l�́M�EY�2����0��"&���<t�z.NWtP5���%��e��ĶR�q���m�z�Oڭ�X����a�HB�T�(���0��i/$rg�J�>��&����}2�3G�^���������F�A䤽���Ҏk�;����K��'�p�h#���\��i�8�&0y��
�5Y�{/�l���Eoz&�`���_^Ƽh�췞��������������m��*m�-���RV���tS�}���[�A�_��z����T����Q)���)�8�7��@K	-y���-�́K�9��vqD��A!K(��݈�UЌ�.
��Yu����.�=�� �a�R�qs�8�l\���9�~�c��?"���1G��[��x�1��{%s�=X��X�����9�;���'��e\�4방bo�w����V�t�$��o]_i`]T��v4�~�����g��c?tR@$��'��?�
�<&R��5M�����X�����q�����Z�,.���`�dg%ͣ׬u��&�	���=$M��Ps*0���\<_��Mh
B��Q�_1�L���/i���j��?i;�h��UG�~���t�����.�P�����k=���$��V��6��WoW��=�����
o�H�NW	�aC&z�f��p"�6��(w�SU�G"Z�]�U'w��+���kq�``� ӏH�$�!���ò*��,��g?pD���z'���-�I�z�7�� �iY�$��~���ٲ�T�!@Mi���ɡ@�>0y9�4Ȣ	>S|��O����o"e�&�q��b�r�݉���V�Cu*�,��o��r��@��aHoU:4��Sp���R����B0�/�)��`���o
dm��1E�7��6��̵�x
���`N�_hd�ƴ�N_�] ��o^�T̈́���~_�!�����������m*� k5�%�L7}U�Lp]<�B��D}X�ħ����G�l���O����Q��_�ɂ��m�Y� ��ܪf}�C�@�!��m���o�h�6�lhW�Z�Av���XlxVHYEB    fa00    1e20u㤇{�]<z�Wp��d.��P<�-�*Ǔ�;Jz[���	.�+�Z�\�C9��lY7@�A�PyS����[�e{�t���/��T�{�+��7�;�@��i�%��4I���5��!��
����x�TF��m?R�����5��GũΪ5��Z\�������1�����m�M����N_��*?�ޖA��1#H+��v,�����Y=�tp�Ƽ�k��
"��@��l��o���ٯ
s
�zۑpX_l��9��`R�g+*G�z�g=Mv=���;�8Qx��2�XZ6�%��.~h�5կX��f��"ɉ���@C�.�Ԫ[�gk�����BĮxF-��>�G�jKKw`�G��Q�$=�v����s�ẹvT���$7�� j�x�Z#h��.�Ԉٙ0^k�H�lZ�h��.�Fz�C[D��ZUd�뺢q(�uؿ+������I:�P�z�b�]z�!^%}4F!��1�mX	��,���Ļ�k2%��Bi�/���79���"���O� ~��"E��M�B@�NC����b�E�s�lM��;�v�F(�Iai�t�} �~��"������������O)�s����5�K!�CRB�o�d��`&p�<�{nXT~�b?�+`����-�S�����0��1|O" }k��j��m�nD9��ѽ�>�U�h��a's�gČ�8#��hO"�k�Y�cb��D���%NS����@h�b7���S�W43�%(#m�K��K�TQ�q��cN�?�`U9�8ۦ��9[x�wJ����I��l8����Jz��B9؜��
�J�'?�u�r�{ޏk�j����}�K�����Tʝ��[;��A:ȽϜ�=&����@Ȭ�)k����#;u���O 7~��׃���¶�����j��'Lt˻ϸ���)IYTևN!���`u���<޺�o3�ê�{��-���$��C�����LzCG$���$����Q���f0_>f���c
�Q)1�HN��x�Y�]3	[G�g$P~h98C	
�X�CX�8�q�XP��vT-N��J�F�q'��|��9�Rs.�dK�%e���~�)�;3���1h��T@�ﾞ��n��m�{� ��G��C�)�� _�Gט��ȸb��Q%p�[%q30�bu�#^C�4Ͷw�U%������ߵ�t�9�D�`�������S_otD!k�d�^�n���F��, ��GN���Uy~,aXe��|�xA��L�$�
��4i�}ٱd;��P�K�A#�!��ĩg��>���Pa/{G["�(����r�`���L3�������n��؊��(%3eWpѴ������G}͉��̄��=��h�h\:&(*Z2<�i�j�ø8�ι�9f��_g܇y-�$�� y,0�^�85ݠnM	�H���Z\kæ����۝��������浩�YK�S��m5{ �	���oZh��A�'V�iI1�g�3����a{z������p����ۀ2��J�����8	��ī,�fCCpU�V��0�'���v޼T�g*�{�3�'����bק������9����+^�wy���7�wQp���4Og��^��A�L�+�?�X�� IU�-��{�6������822�Q>b�)��@C��nKE��qQX-qR�=��ڨ4����qR�^輷���JB�\G^�qnZGR���BL<�AzP8(h,�� x�'Z^{G�C,������mKd7>�v<T���%w�2����n������dJt��x�� 6QE8�P��n;��8I�ɴ�ڕ'(*|��^�i��R��p����c�U⢚�ڿU��j�xw�ԇ�Vd�A3,�[�Izd�4i|�����b�Po����u�'w��Ӏ�;�0�,z��u�lh	��b4/s�� Z3���)#U��s�Bg���G ��x�Ty���K�+�L����r ���5<��)m��He�ؽ��ub�TFu
�r;v~Ty�tf��
�e�Cͻ��8QU��56^�h��4�X�!�0B���5ݚ�v��η�ld��ޤ�廯/�����^f���w�z�8�CR�wl�}���mۖ�mv��'	%趃ɿ���<)�Q��ӎ���E�G�F�~�Ky���H	G�y��My
��b�0'�j�O����=�� rԪ��}��F�`��B��hG��C�"����W%*ך���w��1�C��;x��/3�__5�!R<��%b̡tF��DL�'�ٙ7�E�z�!F���MwP4�u$�е��=m���v����L]��Ƣ�m���ou�zǌ��㹻)�����Um�/���I-AmC�Ƌ�,]%�)�`��X�smǡ�Z�,Kx</�B�$�˖�~�H��T����:TJ^;jN�bO �����59��n��èU�����]��HzI!���&���
/��*�u��7���QW¨�Y_<�?^\�y����]��x��-B��>��O�Ix�<��l��"A��*
%���}��/�+1�̫�/��r���=F�j�p�s2ۈ':��I�|�L!3$|�#L''�i��'��b�.�|?o���:�ōJ�������6c�o�Ä�׼��B=L)H���k ZʆT��lx�l�7(�p#�U��q#�-?P����^څ�zB�I%tO}O�<��z���IZ��2Ѡ{H
�%�DT���"� �x��/�屲Yg��*�W��䂉#Lj�=��}N����V��}]�l�y��d&���˜�m��f����-��W��)!�C�|Uбo��rXw�R�b&e�#�	ϰt��ѹ:�z��nb0n%ϐ�e�+N�-����]i�߉�9��p���|���.x�؛K����)W��#g�:���nR�!Wn!L�a��F��-w/� ��$�=�(�3��`�n������aR���A7ll���p�\e�����c�6A��/<<���P�?ajJ�1�-�Mo`c�UTCn~��r@�i�y����D��X��r��[�uR���(����ߥ��;#�w��um��9Q��������sy�S��j��X�5K�W�H�,��B9�'%���F�W�^$5ڹ��?G����J���pk�s��=Ϝ�W�ۧ�qjf"i���\5TG�#*}���� ���N�3�q���P<��^xK�-O�J6�.�_�NtDA�S�-(f�'�<V���ܷ�ZП�h$7}���D��ǃ�"T�l�}hLf���h� ����!��JΛ=������$=����H'J'|�M�op�Fw�d��Ҍ�4r��?����!p�l�F�w�zИ|���LKT�|�i��_�:���'ˆs,�h\�t�^y��{W�L�Y+�]`-sUc��;��qǙp���,*Ϝ�%s]���	5��f����=�{�J��n	NN�2lk�c����gz� �(���<.���!v�JZW�!�Q�����ZH���8�|V���KL��]��� �Ws����Hg���!�����ڄ6�W9�si> �1���rv���n��Ӵ��6"B<f>B���fab��BR$�{lF� x���0���)�7F���*m2�ntՎ�mm�V��e�����J��Q����÷0�s+,%$��ez�<���'�6��h��Ӹ��c$�!H	��}$�M���x�M�JGJ�۠]K����=n����K�jM9���v׎�Uo{�R�j���2s��k�ŧy�o7������Yꐏ�	V��&B�{�O�q�����Eٓ�^lqP1��&_F�$��ME��P��,�]�)�,�?�l�<��0�q��Mz;���X�xo�il��Y'j	?�>���u�p#�[��WS�U}/(�]�w���z����n��S��1d��Μ��6���}~����?�8P�>�M�x ����䗐D��:\e&y³7�J��0��$��-��U�zڭ��?�������aG��ü�p&�	Ng��{k��!jfF�#܁��몡E���xWO���g��<{��M?w����X9�Ͽ���m��Υ���G��-��|�yRK�#��0{Jh�ީ,�z[�,��L�.��y���y�!S�HB$�J��<4�����m*�[R�8s[���ԙa���-��8#�wP�r��"}���GP�9'Ｌ����͛�pF>�Q��X�p�6�:/<P� ���\��%i@(�#�6��j	H-�xRN�;��U�C���*��Q���̥\�	/$w&CW�S/] `�����TΧ7�?
�;hy��t�@��&\=B��r�� XD���v�S)�p�-�M�@�z�`NYވ���?��R�0B̦#��_���*��r	�K���� @���c�/�����y4�Bw�S~��F���"?D[�U�˫{�V�>-�fW*� ~�-�^�k��J��%"{�Y+w>/o_.�)���Kq��B
'ʃ�;���:*N�=WV���_S![�/�j�>x�yՆ�WcsY�� �����!u�_�M�>��J;��5ܳ����S�E	�J�:��eY=���H���h�C���Lȭ����O�wL�	=н���������E_��*�7.P�H��2Y<SD��A��U��x��$L���a\�s��_��Qh�c�Η�"��>�vC`=*����/����#D*��e��4��i�x�Z����v���m���̂�0xS������P3�dL�kHo����Άv���N9m_£��-�A�Ƨ����nL�k��v�F�Kj�F�t�*�K7W�0l�6>�o+�J̗c�g�����O�l�-�Y�e� A����ʩ�� 3;���א�/��C��D��h���1��T�P�Ƨ�O
O����G����l}�pzJc����������4{ir�M[�����g����by	r��s�Z��}��1{�<�0���j�{�n����K��!�槐�7�����x桞 �Ó���A	z�++�B�7�Ƒqƾ^��m�*�F7��꓍������~H�)���,!��
+���zS�o��e��p���˰�S�����d��A��L�hK�g���� {i�X�Yؔ+��~���v�XG����5�|��(q;2��١z!��B�6��iħw2��գ��]����xG>\�U[���i��ln�]�����;@�2��i6��/1����!��Bf�������6xo�c��H���e4�Т �\i`κ�X&�J9m�t�tP>�nh���g�Č�U��N&���������R�O��?Rǽ=�|a��*la��ۜ&wHᾹ7~56In4gS?�M,�W�xYd{�N��]|�ݥ"n�fE�|{�ep9a�]#�q]�����+PB� 1^�`��F�+��s'�7�9���A����V��ZiI�s�C�*�-�v��j��΄8�\��|��t���Mc�������@6��F��vI+�rH�/�7B��_t�����g�Y��,$�F�)Rlu�e������q;����ks���,���~y��abW���Ӭ���V%��H3/B�
��F��jc�pW�?%-��j@b��uX�󻏞K��\&Uk"d��)!>�P�Z�I6&�V'A�&�����`{;�^�8%#��kr�t*4��[wbh%u2!f���B^��i�SGF(���Q�%��zM�^�	��M�q��>�����//u�����qSǵ�khf�5*�9F���d�e�A�s�,�ыIӳ/"�Z�>=R ��&�}��+ڣ�U�]��c��ψ�'���ҥ�L-$��j'��/��R�G��B�|�l̤%��޻��Pi�{P��;�eT
.���vQl�1{��8e#���h���V�Mr��R�R���?��E��d�ڥ�c�6��c�r���&\��޿So�)�$ߔ�7<�B�`��i���j��t�А�AB6��=JyQ��YSl��i6���,��G͵Rj����	�g�F��;<H���~�W��#u$i�v�B��Km~c).[�-Q̇�����$��� ��:e��7�n^�Y��]�Ǉ��ᚩ$�_��V'�>�'���2 #���èxr�X�ܬ��xl���	�ͭ��Ez��r�A�Q��f �|�®��v��0�����ѡ�vnj*)���\��Ԓ5�$	��2��:�:#{�������&$����d)Q�^�n�Y;�p��W1��D��~M�m�4��XPhȾ��(t�XR�hZsJw�v�\�b���<��-W��x(�q�_��,>'���Uw|Ш����B���[a3$b�I�j7%zy��C�%-� �K�A�@�W�KP��@=t��/A6>
!B�wM���ﺰX+�?P�uw�i�w{׍�͌�5h�G��Fƚ��'�WN�����i7}�N6��qe0Y9[W%���R�)��0XI�BY���7�k�s�C|��&Y�{�
��G��Y���IU?ťC���H�����E�������]|�2;��7�W纃Q}̀�������G����>�2Qj'�h6���
y�u�+��qQ0����Ȕ2'G���D��W��Ǵ��F���` w� ��}ѫ��ʸ��qӴ�h=�_��=X���8�q�!C������~%��X%�sΫt���!R�k��d���q ��|��B��A�eơ�Vg�Dm9�4)g�O����:�FO �h\ڠ�ݜ`��մ�[�[>���i
���Hy�YJ���
�aCq���Mڏ��T`���R���w�U��	EsK�6��^�_�eބ��_��ao�m+Z�A����+��}�)4Y������G��;4Q�4�(���AH�Y+���휇5����mP�k��-��kQ���@[�َ�����Z��A�{�g�xJ�v�F`�`�F ��#��1j���Y
�٠S��qQ%��	�~��lJŨ�d�/;�X��Q<c����Z�_��n��'��	����/ܦ���#_5� 5�4]h,*I�	�R��'O�(c�d�W��`�����KZ#/-O�Ɖ���<zos�nc�n�k��\�Q��]�fɂ��$d>&__��Ac�h?�H⯐)�K���j�97�� ��$��|~UmT i~����5 EMk���E7B<�4��i_�t��#Q>W%�̿fJ Ús�I͊qlϼ��+�hywr ɧ����y��E�p����Hd�
�!�3�"����/���	daH��Z��\N� ���H�}�/�6��cAoX���"��X��y6H#����b�}�r�� ]�]x�s�r���}���:u�L��c��r�frb/#'-.#��:�Bo"&���|��	�O���N��r4"������P9����xL9w�6P��������G�_�Ps4I�$v���.���!G ��χ���C��8K�7�������'�zx����zj^ ���.%$����@�2�+r�D7��L��-��4H4��8��k�r� 4D����U���B����
}A\��(E���8�5�"�A��5\��XlxVHYEB    fa00    1e50�av�T���tՋ��f|�V����Y�1�F ����*��]
I�Є�˝��_��)8"ܶ��y'���%�ec>,���i���҇j�6"Ѵ�p{��L�'O�,�/�j�5`���j�:h�^}Q}[E�	~�9��"��Ψ�X�t�U�J����g;�����gv�.�華�I�ɒo���3��ټ�4���mz��.�;���I��-��=m0?�X�l�g�8�Q�����*�@�M4G}5Se��2��7�n=W�Z���t�i����f�����ز��-�L�VL�m�e��2��9�(�S��<m��.�J��(�E6h9(�Nk_��Ax	��&�>}����� ů+�=�����;��=K�X��;���yO;�b�	� R����)�4�	_4O&$z���n���.�g���1E��(9�\r2����F�Ѱ�R�` �F� �bG}�"�����aE�*b�m�r��/�,b�vV^R���[j�hyp��%��w�Ms�|�f����	mA�|%�# w����
Ipj|	��؇�y\��&�?�g8���ovOg' ��eV��B����r����Uَ��(��='�@�X�	�B荈�2<u�љ��F��kҴ2��z�J�?�A$@����f�P���2�49W:
�\��!���$���=[��"̴��*x��ƾ��z�}�Q�}k;���K����Gכ`��&��w�_��O5H9����⵫�U	�X�:�-�:���Xx���,�y���N��h�P��-�.v!e�ɷ����<t�`�'�>K�8Cyg�:Ȝb��zB(�k���<���y�x���r�r"���1��< q�~��J?��#"Z%�B����4)�,�<
j�Xa��qP����ϧl��hxe`�U΃GII�!�W��!�jn�+5�|�NA;��iD�����4�鰯!��ʮ�s|�6dA�Ğ3r3�f�"��qa(���v��ޑ>M*nY�ޮ�A��?DL��K���<�w-	o�e������&<@=5&�ŨEiH��#/�f� �a �3TT��c�X��6s����Ed������U���X.��̱�	�yl
�$C��;v]c�1�oq��8<��A�l�%��x�cX/*Dݯ�(��F(
�0�r(	��ٛ>���a��q�AL|.����B�/�����YV��a�R-2u�& J�����n/]b��ī��t>�M��PBy8ox�����]�;�9�l�ް�S������E7�$yt����Oo�B��_��/e>5�ˡƐ��0ʷA�E=�ȶ�x%~t� �
Z�����r|Rj��5o���
�W�-��^����S��S�9�&����~���^���ۮ������Iv�ݟ����
ۑ��[$\?�,�N��9����bD���o�>�u{�sRtXI��$k�{����5nX�y���o�"y���8�{;���-�]��G�r���1�&XH?[f{���i��������Έ��5�H�UO���f��o��Ir�ʫNti��vGJ����yK��Q�Ec���l�w���p��^�l��X��(�r��,��%�=�l=����}��_������=� XIv3���~�G�84��v��� }_���<!�$���'��HN8s�=��-	j�u�:�N�<C��H-B߱ɚ�T���L:�u�����Ck����҇JO����P?D���|6�0G���P4���W���- ��s�nj^�>r�b�
��j�.j{nS�z�*��`S3֝Fh�ߺ�V��8���粐�$h�m�]�ATt�*��9�W�5� 0L��a��0�%0}��+%��'�L�=�Q ��HT�Ga=� ���!\���8�^�C���׿�n7�n���vRɖ�g��>�꾾�,ʨX:��4nb�1���Il��mA���$�S{�B��OL�$�M6�5���f�g���Uq�/@�20/��9]��o��'ٲ@�m?��3`}jI��+�D� A��@�����ҵ5�4-����7_![5�~�p�q[�2m6����j�L�`Fr�s`�a��2/a�g�~t�]ϳ��
��5��z����9�{)��d��8���C���$iȌ���n%�����8g��ll�t�'x�W)�ycI�R=tF��Ax��{��cůC���.A����o����l���W�}B���t�n.0���8�g����P�R�\*;����:E.�u`��L=+�cYD��qsa����=���1�B��Cf�{��ILS u���,�� 8�x�%H.�"(jz�GGit���d:�y�����)����?_���BrBřW*|�
1���7�M���dI�c�g���z���
�&�L���ᡉ.�S�Cu"{I�kaK�rb�!��V*o�����@�e �-�E�B�C^tH����GJm�qݕ^(Q�A�z��cˑ?m����Tx���z��� [�\-�aI��dqN�N�tK;��o}�����@�����JW��Q��T~�
��^���#,1����4R���X_��(+��oI��ݞ�E���\$ޱ��x�@�?�q��lt�np��'!n^��W+3ubbq���<#��?�qK!��슦c+�B�Ym#L�a���HF� �;Y�P�'^��R���x]b<��H)�'�g��?I�A�m�P�[��3�)a�~�]�}W�L)��Y����1�=�c��h�k|4��+���2�%�7��ncT��3\��!&��1�H_W��qb���8W��6�Q�r�A�������ȺM r�  _�ˍ���b��4 1�V� ��$]0��oH�im/&��fc��3iT��������o��*.�
�_������g��V|�0[���2

#��������b�\Lv�<�Km{YhK@A��gj�@�â�Ѵ�K֧t��g��BM���۴��t�~�M�i>�X�r���^�Y ��n�����j��F��	%�,�m��c՞H�9�a���f���V���̈́t^"�@v��3�����A�8~5��[�n�Yqw\;��M��X"n��E7�C�$�fi"�UGʞˮ��(�g���E��NՈ�͕�쮼ɰ��T-���C����|�9m��X�ۘ��R�{�B��p����,η�/K#[C<�Ċ�p6��q����p	I� a�ĭHr��ԩ�qb(�����UO�O�R,����Z����P#"߈/e���k����B���d&@5\���	��9�(	�\�6��ӊ�m�aRB����rX��h?�}�6�{�=�A��I@������ߔ�!��N���j�b���I�0�
�[�����e�¼�����hbtݟ���]�L�5'+�i�޹}�P���}�rf�Z�s���c�;h�߰k/�����,ȏ�e�h��zvu@��tfXGs�{i9��f�4}�2�I�^zdw�)$rU�٥'�-2�=���E��&L+�ڶç��y?�y�R1�,�t�Ӥ����T��|���Ŕ`�-\PPr����w�4����I�N�D9��n�J(cR�+	nb�$C:�Sap���j3�w��ȹ��a\� q�����w����i�VT�m��^�x����=�s�{��Ȧ���8�%���6v��F����n��qs7����yS�SB"�}񿜐G��_��:d)ap%6����j��۠TE�o���� �d��y����e�@�_�3B��O��ujpe��pW�R��w?�Fw�#酳6�̽�s���e,	u��*�{O���fx�E���q���2W?���f��9������Rv�N��D
u�2/���J��W�z�%`Z��O��p��Zx"�>�(f(���T�1Z�3�ح:�	�"8}}��a�9ʺ���dB�*B�+٭c@�,���W/C�.��q��  /B��`-`�x��ȸ'��f0�9���,�����gF���2�����v�[��ɾ����*�{��R��:}ǃU����t�� ڜ���W���R���UZ~�V?P:K5���ڠWD��j����� +| b�ĬI1J�(���
W�"�ńE�9L���j��O�ӷ����j�9<� �D�R+T�^�t6��Z�-B�3"����(����i�|�j�=�0�!�`��C�&��-�� ��W3Ṙ �kt�Ka�D�>���xF<�<��i�RJ̞�,En��"�״��z/osI�;��:VyJ�x�w1�]��ܾI��;��5�hͭ���q�2r[��H^�Qa3��� �r��� p#15LN�vN?EС[p��۷�� kR>�_��%���6&��vn.����I��q�������!'�}�.�q|&E���R��J5��o
\-6'��8�p2D3t�$��R�%���Ng�g�=���H{�ͅ6vV=Y���p�|,	�Y&�@��;t��s�G��op�W�eu���/�	k�T|+�-����q�r9^�)��8��!z� T���I��S�]tl��5�\��CN�@!{�=������.����V��!���?G�¥���pY�$��uT��ϴ�C �?�c<�٢Y����Q�A���
��tZ�vsX�t�+Q���&@�~r$�;��(N���,H(1~�'��s�E����0�����@�v-�<찵[6#̜��J��e�(��w�pi��0�v\%��E��q'�:P^�(�<qvk������;��񯍁�L
uS}I)$����?�W�~j�&�T`4�}r�l��_OyD��Bwb;��̸ݵR^Uz�c�,>��JEma/�p�bG�P�rEF��/B�Z�'+�3�R(w{S�!�vw!g��i�ɾO=�c�"��4+�E��j9�&�u1�������z]�Ƴ4z(Q~dQ)�u��ff��@���nR#K ��wݙ���BBQ���"Vc�Xi����P�t���qsK٧�ϰ�F,��C^�_�O#	p�1-Fو���/�W�W!�-b��\پ�ïvTa�P�JZA~(0�G$�ocY��P�ֽ�jg��6e��:���F�)�����[��<\W�y����H��rl�ؽQ��D��4���i9o[3-���,��%U?��^�K>�T.��8�5'�v���� ���O6m����m��y��Б����( �,��N�
.�&��L�#8`Pj�;��3��._�C8x�/ a���n�l*�w��]*K7 �GG��G�zC���Y$�5
�Paաu`�b�+��5�{p�
��^01�>3xz�Ax��vm�ۂ��Z��rhD�<�0X��Y0��6`�ut�U�������xb_v��8Ѕ]�2�������z1���t��D��
�R_)U�(O����:$��4�h>D����b�j��.�π�	�Y�I,Z��e��BXª\E�S����1��5��RqSu��O�,T+��n�����$4���`Z]�\�)a=��R0�eE����O^rD <F���yc����V�f�9���U �i.e3��1�NB&�3|��L'zob�R�f�Կ��"�U]���e�^*`���Mu�~�F�H:��~$��Ο>^�5T
ߠk|���-9f,ejӏ�J�'n�}�h��������G'S9��6�����ܜ��b1<�[�F+���^��)#�ɵ�ݤ�}Ih�z��D�bw�Za��r�z��$Y[@��u��5u�� ���4|��D��R*D�v��?{g\��W~V��̧@Oi0��~��Ē����4��,FAZkrh����^y��:�yK���u]mwO�7��Ef��ڳ*��W�+�@����@o��6!ʻ�GҼe�__W�����Z%Ak��o�n�����j�()/�+���������]yAL"�W��tuK=f�|DB8��-&w7�y�O��%�Ҹ���D=���C�yl�U#�5p�i��Ѓjܘ�g�x
C��42�h���TO�
Y�q9_K��%�JF���9�k�8��,k������l)�ƴ3T�BXi_4�(҈]�kҏ4b�u^�Ҷ6ʒ�� �a��[֘���Iw��ʵ��(T��������C������y�[��IT����Tdu����)��q{N �b��? 3�b�Vގ:����|�!� lF"<c� 늞y���%�l��
����"C�A�Gs6�����+����
�q�a�*���.�kL��M�G��|Ef99�H��b����	���үLf���'�ʤ�`y��:�	5�h���VÕ3o�o�f�ʨ�&���`x?H�Ii=s��x�{U����j3���|��4f�}+��U�6h��qs4�]B��W���"^9�R��ٱ���!�d��
�E�� �V˵�)���`c�cs=+�E��,6�C�&���:��}/���JU,,�F���h<c��K��jl6��Vsf &�?�f�$!p�S�΅�#K�:��Z
�&��Ox����*�P�A�*�gv��I��A\Xﶺ�-;��(�M+�k'0p��bգ�q�U��6L�3Ÿ�������x�4t�,�h <uѼ&�cJAS-��i���5f>}�|�Z>����N�6�&*{\�t� 4v�8Ի�r%��OE�Ng��n�	��/_��G?`ȉ���{��RJ���~@VF���v���|0�wF�Z�6!�\u��ا>��Uّ�	6��������L
�R�%<Nd���ȟ>y�f��#%BA7������]M�&����>�5��=��Zi��m[1{���V8@�5$LK|3rj�k�����6)�Dw���H����%�mD>���xe/���D�bo��:!/�(��V"�/di��(Ԓ;fg@�0݌�7�?mrZ���sd]\I�j����a��HP֋���Y	��ta�:��{>B�*H�P�7w$_ٓ:��$�jo�z�X��	7�/�2=���
/0W<@aW�*�����w�%�Bޔ	�|j�s͈(����������B�~pf����)�^�;a��z��A怽�Dg�q�I%���Jt�I�� �.+�3���q���z=3۲�����ܩ��l7���f���/u=9�U��n��A�v%X�Ɯ2!�-;�xC�L(��\ĭ��m��]"�|z�|]�ӵu�iƥ��D��?��K&�?�Ke��K$6�m�B���i�U�?Ν����}��cr�-�h���q�ŕ����@4��8R�f�J��f�G������z�@���0��[w���ǉ�%��W/P��)�@y��X�	�%�(N��Q����Œ�~:v���g������E=f�Id&&5�@��"� �Y��߸��ʬ#W���%��	���T)��<rϗўm�ԋ#QX��յIE���{SM�.����x�8L���166�o4��%�Tڇ�|�D��Ws�Q���p͗�%%N��p��3Nw���ks��M��я�?�	t�\��\)\�N0�d�	��p* �D9�F_�'�J�<���n���p#�-�^|�4P��F��n�I�p�� Ó��1CY�2t^CI��Q�~�\҇}>W�*&��6���&vXlxVHYEB    fa00    1da0�����Lo&�J�
'�+'-��������'�.S�n;��LJz߆� ��عq�Y^y~�\d�~��̇�j�A>2߃�{#�h���͟��9��wP��Ϝ����uپ:�i~UА�f�T+i���6/oag#s�mĉ�֟���J tmI,�$�\�[��<�ܿd8cGҽ�@T%�bx�4��bÙ\�P��>��.�β����n`�����j߿�x�{�w�_li�,M��F�˼����]I9�l�$��gEF������m�#������T7Fl�k�2���M驵�eV���'��B�V�i�$.]Ӳ���HT,�N�o4a⣮_8ez�\��T!�s-�d�J-_񲖚�����j�6j��J۽4�HK����Q�lбwl��{�����1I��U"�)]��!���V��Р�=ѿt��Pg`��i�F^��/��r=K4��w7B�		Wv���xA-���@Z4��U`���3����4�W�<�?��X�7�"�i��Yݜ�q�\EF�0p�>�3q�	�J�W�@2x7B�4���Y��A�CF���T��2�l�����֙I?q��&�p�]b�O������?_�]����>Jj�/�EN\`�OT��{�"�;���wѮ���/��ziog$�x�_Q��K5 9�z>D/%!k�4@��+T ��8����mV�R )�S$��R���(�f�X�.v}2���^ސDCU�y@?)ة��j 4�tD�����yУ�|8��bA{�ɼxX :il��F��������p��9+�3�]r����E���;���CJ��`F�K��������3c�E��	�Z���:l:ɽ��i�g�^T����J�F������yZ�vO˒b�!�qar��~��O<����x�6>�L��E�?M2��;����3���d7���W�1����VF�����|��/l��� �o��ۨú3u�*�~k�-���jz��	If����|]b:�b��F!�Yo�c�AC�EwЎ�Q���,5S~�|h-�+f��;�V B�;i����r0�"z��o,%�L+ޕI � Z���z��%��h6���a���­�W)��;Z��vG�0$���4"�,�͉A.��C���`h��U�4(B�s�=|�Z�(~^\NN�}�U�|��h�RU�Ø���/o�����lQ�7P�|����4iM`�3��]A�o�8w�@���p-�_���ā���UzA�
̻��Fi*�K�9=�@>{#�?�?���+����k�d����y��<bY=b-��AՐ�gґ^��y����zkLV��s�!�ƞuЇnt'p�����"S��E��~���+�1������Q��sm� ����e������*K���l&�1H��5��@(���!V�=$�ZR\�W'�#������ٸ�2t����t5���I�%B�] �q�϶�o�l��к�wiV��Im�R�!��%H#2s��`�-��F�zC@�Q��X����,���q*z|&Bq�k���"Q�Z豶������c��o��טx+m>�@Ϭq�+�����s�X���ϗy��H�,qO�&����53J~М�H�!c&(&�D�%��>�T������xՕRA���)v#�|��K�t:a�_M����AZ�엒-��z��4�%q��1\m��m5=|�=�/Z�n_H�O���RwD����Nq���̛�@<c�C��^�ОͶE��Aj��!~�^�U��ϰ��<���2��*��d_�o���M�(��+.���M�nD�*h(�9��K� �8W3�De?����yCPS�
T�{!�����S�����(�_�ŕ�k����%}#��EðĦqh����-\tc_����M/�J5��(�����/�����c	���4N��u��o�}�*��ll�� D|�;��wbi��ַǤ�2�G��(��I�nӕ��4��Nv�X�Ӕ��a�%�`�:�)��}�,�� l^h�;�Fq�����g�h,Oy�̖�"Kx�a��OX:a
`"|C��:��m���2/������Ƞ���ѷ�2��O��9V��-BQE�h�3E:I@|�H���*>tb���� �2�T����[�ve�S�������o%T�Ut.�zt%�ոb@������M��'��]��U�o-`��#�)��/!+��0H�zu�#-��:��p��;uO:��Ygx�$+^I?kw���J׵�kO�俤~�)���z$�4ٲ��%�h�Л�Oy�$��FTZ<����d��h���o��*Thl�D!uO]4�_��l"�6Ķ	�.!��1U�}
t߁�o�b�$O@V��3w4Fw���)H�$X<��W̳]i}
8#�pp��^�PQ ���������,%����S?	j 齙^\���AUn���
]j��@R�w���� �=���F]˂�}Q����*����7}����s��M���N.���>j�c�)"�-�Ly�#PW����+5�2�^X��|�� ���G����GC)^Cts�O�xI��'���5�Q��5�VI�J�ţ'95��YBؿ�=#���T�s�}�[:�Ҫ�wz\j�@�A��)�;׃��E罠��z�O}���+���L�;�b��=����d���H���GP�a"��*�/-9�,�HS3uٸ�%mC��x��	5ǾmxM�
ie�6
LkO���]ǰ�Uk	\�"��N�Y��2Y|�D���'A��iv��Ӷ�tO���
n�5qK5�� ��ôsD~W��م�I��ً�!��Et��xҩ�����O$�wȂ��џ��u����A��_��7��I[.ʀ�!�g���v�]�I�S�UH���y}&��V�_ܬJD��p�r�z3"� �_�"�W=gTc�`�L�|U]v�������������IͰU//�>�Dq̺��(�1�+%���晢kt���ߡ����o�,҅����%1����6���ǣY���*յ��ֽ�o`�������X�8����Pג���bj3����fi-N޸��AQ�yR�AT�l&�9睓��=�*t�X�zC2(r͙Vާ��yjNn?��\kJ������.�[hc��v��+��q��'"�%��a�����V�2y֪�|��r|��7�h�>�#�̗	�d޶�b9[�~�Jx��hy��|������$�r����͆,���݈���y]̷�N��
�˝F��@�U���������if���"Q1�b�[�\�;L��0��h�V+j�[p1���{�Fd��vz�X�������u6M����ɣ�?�$�o��#��L�����g}\���ʷ����U��?�C���e��f����S�_N󡁎�怯=r���=��H���h�_Q��P�|`i;a_l,�g�e�z��Ƌ���4��}tIͮ����n���y��Co��ٖ�R�i!탅���MS%e�˶t���u�7�Fc@�lf
-PMUu-W�Л� �BM�c�s�����Qq�B�Ͳ#�͍��������E�z���yp�kK2,M�C/��݆��"�l�;����.��~a`�#?fZ����0��2H40�C���~��\�K�s����.�UP�Nyc��ĞU�9pدX���?��V*:�II�c�#p'����C�<I-�̸���^��s�{7��"Z �fi��&C��b
�nH~�;%Z���e�e���������jީ(�8��0��\�?�?;l�xc�
���J��{�]g�����U縚�TMX��Z����(`W�I �%�|+�r�Qb1�����W
�Ra�uͅC�ݟ�+b�f��L��� Ej�B����-��G���$d�}A��x�r�I^����6�fLr!���:H�xH �뭢}����.:��Y��V(�����JAٮX��� ��gʘO_&��G3���K�雷�^�`����|U����ȱF�3*��(�_�*���|P!��&=¡��kF�Wϑ���[���~�D�R��Sb���dre®X;I1x)(6�\��4��a�C;��O���'6�/ J1Ro�8	�9� `����$�e�)Xg�W���2�X�8����_�L�������ܔ"!���(Ts�u"�g@{
��ZD��"��f�"�3ҪMOתĤ�f�����ܽ����G��Lחi,�	=`�|"�V������r�}�ǂ�.��9v��n�g&͑}���c��K]��5eD���I4�1r���<8	��MԵ�?��o�}�hX�73�}��n�弤Z_w�>�(��~= ��L��w�f4�G�����1��ЮQ�2�Y��U5�9��fN�d��lFί؁�+��M�`IE��:<�?���U�t,��a���/�w:���?��?����~m����6�����" �4� &��j����C� P��_!e�G�c�v"�=�ވ�_%	4dS�v$�ky��������chk.�ȵN��qwVm��1��2W5$� AI?�e��i�w&l�6[����:ɉ����ߘ��	փ��;t�5����RWXMq�[�������7�c��c>�S�ˢo���L�Oc����+J93�X�?�z'K��ǂ,.{��G[)b�f�'�FE�h������|�)Zv^��h�f;�?Ciy'�����z�-�4�|���@f�����TՔk 4Eb�����6��0���sꢭ��j�z���&�6,�<zj>�jW�B8̳��g�p�#r���5#��=��c(���,���3�@���k�S����HeLWFG�Z�T�A�j�/�ky��k���Ӳ��0v��G�ȷ�N��r�پJX�l�Eb.����5_hFɵ�t�tC��(��=^�rd����%⦑�U(y�U	+'�OP�a�C����{�'�S�<�K�;wO�qU���OSv�k�}�e3��f��#b�p4��f����c���ݮ���@$;�Ҕb�C��RJ���Tv�� M�c�y R�oˉ�2�}��+�ı��K�A���U���<�X.���=>Z�9)VB������	��������"�"��*?^<�v�X���1��&�.�ص%��T�m+�^SWK����s���a�J68�d�`�i�{�񕾴���j�9��H6��Pq������x�˚t}g괃$�OL����0`�s�o�"t��;�6N[���g�\�8�^LI��T�*Df�ڗ�ɒ����O�8r��]ۨ�u٦ѹx��02�^�iAU�G�0
���5����	z��z�f{p���*x;�-�{�Ͽ��/@�z���Z����,0�2 Z3Xg"Q=H�*��7/�ޑT�x2'�}
߈�Um�Yk��dZ؎��������d�:�}�R��,��<P�̻ � �9�^jtE�5DV�ld7�暼�&��e(R�:�8��D4�g���M�h�S�	�w%lVgDUOQ
|S�9�!�����v`M���D}�E�D�-��ٷ�O����Zyc�C	e�Tr{j���QG�x�c�Ө"���^h������-g�2��}fx}a�<S�N�U�7a͕	b��K�	�=��[X���0��~Rgz7"7ў�%�=wJ)y��p�7�Ir�԰u�������1¥]A�I��PO/53��v��x#�6V0��� f
H0k���<��_�,Qhe����](����{%��M[ON*S�c����}�	A��Lx�T�¯	r<	����u!�Q�����'c�pô��.T��D�����x�O8� h�Ul�?M��ci5du�1ÔAUw�Q��q*�O�V���`-�����Ep�)H%j귥��gj���Z*���U��`ؓ��.L��yɷS$	6�:W4䅤����~(,M�fd����V(ϕz����p,�ͤ�aq	B����pE0M������~O�F?�(�
E��I-̕c�ޮ��ܸ�j8��rv�5Ǔ�"�\�j��U�cd}��F�c �s(qy�T`0%��B���|)�VzE.���H�p)jFG�t5��qx��ǻ.�%���ur#j�:�_;��mZ��⯱��}��N�(��e����z�L������qz\8��Q$]���39k��cA��_�p����Y�i}ꌷ�a��,6Ӱ-PPS�o��>Ax�Sp��8��K`��&G���M�n��
ѵ,�����P�̫2�J�qUr@��޴��Ux6l���3;��TZ����G$�� �h;�Nb\Ypo��,2�H�^a޹��r}�\.��f�4l�Ő�Gn���.r5��caݲ�TNG�	Fys�۶����␎M7i��:)Q^�-rd�8� �b`�\/�Jf�p3l� |�����4P�5�����)��ow,����̤p�m���X@6*��敘�K�2t��E@ve�n�"w���"�^�!
9�x|R�7}��h�3��R�ln��E1�R"F��ͽ7�O+��C�T����6����T�ρz꫙��M��Ӎ���Nl��Ż*f��_��iR��y�3Vy�}(g$��p�VE�a�l��zb2���#�	�󫬓�pOY�߳ �9�jxB�����༳�#U���L�7�1s�Qa	\q�P�aG��|&��b��͉�Kȴ�IғOF�c_��x:�x3���34�PA�ك�O{�ȍ�L�s���b�:�Y�`�za��K|}/�@�`m�l�.UC��L����-�����3x��)��}�^Ȣ��S��4����n˴9��E����ݣ��������I�+I������{|�:�,�v�m�cCgu]O"-'Z9:a�����K��f�-8�<���P�Ұm��㐑���Ǟ_l	���U�5u�{3'���ٻ{u+�'�Z^�|�GB����a°�&_y�V�Ϭ�C�Y���Z%Z�G˹!�񡀐��V�a}�pM�QP�j����R�:�O�ꌹ~*�����q�$&�JE������Ʋ���dt�l�e�h���Ƭ��rϰ��E��ԶGG��_&@j��H�A69�>~�#^�#-+'�S�NyB���߄?p��3���5L*�x`���Ob��#�fZ\K��N��9ӗ��4g�Q��Ի%�⇞�$�gc��8N@�%z����3nW�A����!�H��$#�c�jt4`�]�����d�s	rN؎;���),(�s,����nt�����zɮ�'��!"��~���tBK;�o��SC�|1���i��(�l��M^��F���&��!�
�/�vK$��%�|5nuߺ����l�m3b�"�*�;'�]���Ŵ���X.�,R��d���|��#��ڧ���ծ��c6n�eW��%e~��33��?�R�Ϧm�bh�s�85�v��A��&�T��RC�V��C	���r�K����XlxVHYEB    f314    1b50����ݙ�%PC͎�H�� �6�f3��/������4E�h�E���]B���ˈ��O>V���IdB���r�^g�˨�H5A��%9���:��^:����N�:5n%':ے�6�&]���Z�@���p�lr��P��JM���<��+���k3�l�.\i��$�1��_��4�V��Ʌ_t�7*�-]������
�:������R2�H�� �Q�_"���%G��,��0R�x7����p�C��&� :�^,�޻d�qI%~6��$�����{��rcM��:�Jd"��]�cKC�>�T��l�+\�j�L���hK�����Ѡ�� ӏ�n��8���d[o	���O�Ǯ n��3N�C��+��"���"��[b�dD��r�{u�O�R6�u�'�S,¸_�d�Ĵ3Q�Y�[?E"RԽ� ��/hu�q.���GD���2R���X}�i���;����x�U���[j����ӕ� A��qG&d��N�,��ܢ���J��'��U|��>w�#I�L�L��nK=֘A��%�%�>�Z�L�Ȅ�n/�S�CHnH�"��)�AeW������/�玻�=�[?�����H�v[��,\v���ֿ��7ղ���r
��16< ?<�;L�7��[Tw�/�:A^��y�lWZ̩���J����w�	ˠ815�	�A��=��"S̏�PK$#��Q�ݒ1Y0����aXn�};�7�p�9���칭�,Aɢ��<vmG����ȡsg[h�k튾z@M��t��YR���|�����I�\�(��b9��4����fy`V ����F��HT?b�Su�ZG��d�I�L�Q���T$���7Z�\��^�XFJ;�볩���na���(��v[ꐸc4i��H�J�7�j��rG�*���3�ќ1��C�I�R�J-�Eֽ�٣����4d]�a���k����O
���(�%������VBc�w؋��x��X����r���z�:��5� �W��h����<�͡c'�:8N��L$�$8�qL;6�[i8.�����T��я}|�̿�y��+	��c[��:��W����5U���Ѓ�2�t��=��C_r-����U�VO����.��tjbo+Iˆ@AL�4�A+9Čg�SdIW�[q�F�`���@��Mj`x��Qn�X|؛bW~�VYf��>X}������5=f�j
k��9¸�Z����A�=v�U�ODA��X�[^WΕG�k�+�j�𠕐���&��*C ����
|u&��}E^� � آ��ư� �K�l}PqKq�%X�ۦҷ�!z �l��KB��*�N��U��#ԩ��ۖ�^�����%���ց�����q��hR�2$��!���g�����j�hO��KdeZ�5��$M��z���ow��Z��uE A>e��-Q�L��YLqG�Lծ>�+�;����z`Xg���v��cG̒��\/'n������hQjº��P,����Y����e��)G'w�����7��i�-dTIS}pD�O~��8R1d����句>��]6[`u�'����*-�"'�������X�x���Y��GJ���ӡ�M5s��KwD�;M�"���n�*�����s��2�A#���2�� ��+�����iU-Nv���W���p�-(��p{�j�gz��d��/��	O��Ge���=Cu�.6{'8v�M���[2Ѝ�l���h�*�F�j��3B�=��]�F���D���aZ�ա�����E��&��|v1���/6��̝V�I��/����H/Q�0,#�T��!��0��S2�̶�I�O�d�g����N��*�f! F&W�L�=��i�=�MCp�:0��1'����q��t�mc@�᠐��_v����[L��X���ld0�H�^撈�E��ߞ�}����.�0]��(1wS�g	 ����oW��s7C/��f�"68) �!_w��s�3��HP]Mu��N�?� ~�l^��E+s T-D����]mMZ�t�2l�p���j�[��
#����ɉ2~S�����Z�b�� �@�J���]\`ᖞ�������D���E��T4���y���x�F c��|{5��_�L;o�̢�)p��?(�}��ڞ��m��I�k�������;���� ���6����4���Z���x�w��qt�aܙ��e~�f; ��#L�.�Y&9q;t8�[�ܮ��A3M�%�PЬƞ��ü(j�����,�6q��"��݀���:S��t>����4?��5��+���2A�Y���up���~[�X�j�Oۀ�~�4�u�,=��T�4��
^��>���q�X�	��c+���Q�� <FB\`�U�����#w�mc��ݙ��E@SKK��O� �}��g�@l�<���ݟ���[X�k�w�D ajD�ؚ���f[7��v�W-i:���K�2�k���H�wG
TR��c��o@���漣Z�&������"��o��[a�B�<��()&�k�����)4%}f|���j�hc^WE<Q�D�,\I�;�-����ݮ�yp/=1S}ѰglOR9Z���M&����(��o�������|�k�����?����.�C�}�Z.a[�P��i'��k�m%�5z��Uhn��8ڤuC��c$�;V��I�-��(Z��0�sQ��d�t�`B�+ƆHJ8�H�\0�������C*�1)�u@6�=��?ŋQp|+qו=�:(�G^J�����ڬ�bPcal�y�mdN0���ܦ~ נ_v�	z��-��J��'�?j.�W�IXl��<��4��4@c	� ��"s�2Z�c�~z�� @��0�����Z[�1Yn��ه|;O��\��ϳ�����9���
l/��	�%���R4�X䘽�I�'*� +��v>:Kf�UV��w��������{�H��1ځ��*�E���d@�����5ͮ��E�t��"��2Iu�|Dg�����b[���I��P.��J_������Y1e��lr;�W%��j�����-�*��YRx��ԙݮ��K?Շ� �=�Bj�P�Y�E�vb)��d9P�<���]S��\�ԟ�.�����UY2�b�R��rZOO��%g,�_D�A��9����kW��p�Q�B���ǜ�C#���g��
���n�Be7���9E���{�hA�����c��FA?@�d��@|�R�]1�	�ꂝ��&��X�u���º�Ks�����:&ꐜ:��V�t���T4 K�����W!T�cT:�v�!�wwC�U\��R��\T��78���H"�1�&�ٛ���1�EW$Q-���jʍl�>�M�.���m�h��ֿb��U�㮓6��gk]�ёJ�u�1&�#��(1B�t��+*� G!N���w��*e�ׅut=��F�h�*��M�.�s_�IK�\��V����F%��4�c�ʇ���_~gT�C/K83�{s���3��^�J1g��l�	uVSza�d��Ogʖ2�n��l�S�b�n�瞳��d6�:6=W������1��g�D�c���j��(3s#���mK�yK  b�+��oZ�K���]��"d�4?"�ҽA�+�9���4�ͫ��3t
��Y'Thtk��Rp������fU-]�C�H@�)�jw<�CFu�2�\��y1w��yq6��]��ob�NF�bw	g�Gd�C��Ct*���y�Zm<�3��[��ְY��"���CGme�+��4B��WE޷�3�ن�P�#��0z� ޗ&�\�H�_�e��e�\-��It1\˻���S3�$0S\"@�����%�QrN�6�&���o�������c��(����?^/�f���HzP�
���@`fw�Rv�t����`���)p��?�f��?A�S}L��Sgda퐦����J;#�4�M��=B_}Pf=f���^�=u;���@6�s�{����`#��e߾kxB`%�p��E�H LɚD��_F3t�t�|�v$���NR��$y���Ե�8-�ܻyá<��S�P���a�;7ϫ�xLPG4O@�JW���
�:y�Q�k���$�0�-b�,ꢖ��78������N���B[8�����V�O�6�WĨ�5΄��=�)�G�n�3��;��k@D�F h\B��/���dk�=��{��"�ˮ�{P���ϱ��(���&�ȶ�Ę�~������.��1�F����Ε�~��K��sQ�ה�țY��J�}�Pp�D\�fM� �vE��Z��)0�2p���~�*�,H��-U��w��%���Xj����
�-n��f���lm�T� 3ʐ5���2�J���OT�{:�I����^52;@�
���E�������&H RW�� %��iU�l��QxRr��"o��h\��os-F�����O纮�q�j^(�Y�o��{6,�mp߶y�%1���ђ6�v	���F�-k����Z@`xoN�v;S8k��/ƨp^
#s�eͯha�	���r���s��'0g�_yԟ�d���r��8bO�'��I��6*8\n+����@L���c�M7�x�/�.d�fV[�^&3(�p�x�,&`�HcP�0��@<��n�k���k���I39�6%��>�͠B�y+���F�Rp�d2��5���������a��m�,�y�&惴3�+����}�q��~�x���2/� %���eX�3�=/eRS��B�g�V;�dr��r���"H�AUq1�]|ǧk' F���Y�g�� ��	�L�˧	hE�����H��&V�l}��5h����W�2��V.Ԍ��1�e���܍���}1��V���z�7,���Rx��	���p�A�`�١��7S�Ci�y�����(���V$`&a�?���8�����C��7�P�|�Y�
2	���(paըx05����=3tDd|��<�m��^��v�	�b��OY��?�Dn��Y��X�E� ��3��>�U~���M�F�y�we&+�a�n1�f�oP�)�͙ܶ"RvڒG��{��iZ��؈V��F�;�X�X��+�J�p��v�O�����"NF�g�\��Q~�����9�����/�t��r�|�I�57��[�!lfb�J������P�|�PAj���{8���%6(C�0�`��pJ�[r��A������(�U�@�+�Y㾏�l���@g���-D�V���@Y��~�|л����D�OU�I��P��5���@.KW/����/�w͛ȸ(
cC�>r�.ڪ	,��^i���Dӫ}s8�� �%=�����|��	�$4�k>ʉk'�1��8M8��!���0M�D�Uߖ�IXƊ�M.G�?,��l7�[��FnWR/�[HG�u�[^(�)�}�x�><+��|��6^HSP����C=˭ee����T>�;^z�T��+&M��c�W�z��\KF�{�gO��K���hb��T	T��坰B����Y��^�A��}P*�8��mE�?q�9�&���{�'I�;�ǻ��ѱO�p � �y((J�hY�~����������M�ð�S��T�oj	tYJ�^mx���\���D�[Od�"i�!X�q��BQme�(�c^�P���\vw�N��F�������׫��*�h���`�ܑ\}�VI��4JE=
@���R���?��������P��b��O�vQ��������i�7�\rё��(���Y�mX�ҙ�� �U�S8z�����"�n�C��l��m�l��A�d�I-Wؑ�-��ݡ%F�����2x��+����]śoK�1���)��U2�jV�C�����xuͰ�H�^m��zt�+��c1c�`�*�v�]���5��)�R�p�Q���u��<� R��z�DL�
�.Ԯ��\=		�������J¢j� VZB͹��2�'�D�Z'��z)�!���?�E�`r����>����h�Va��t&7}, �
�������8�%+��v��&,
���I��Ś�ҝU��_��>MY/8�6;�.��cU���7�<�-+@e�-ω�
�$��C�XѷS��~ɯ���x�`���Z�%U�V��LYc��K�x*Aj�	�wK}>},�6V�2hx^�Ǒ�w|�I�o�T�(��pK��#�C��
�l��1�I˨ �-d���8isY�^��tz���_�R��F*�p��0�[B�j��jh�^(�#ǦJI�hA#�)5�F>'���ȋ%�^�c�L�ty�H`�/ q�.�_�hQ�RCE<�-"�2
T*'�c��8b�~�o�H7�[��,O��k6d������E�6]�]Y|�Sþ*"���o�� ����_R��`�!�#����|�4[.�g�����疞8tid>1��OJD@-�߷�|����@� {�O��ň�T�^��i>���K=����/b���W�g��}Em wa*�$]5�'n7|R��f0kcR��d���̥��M��Z�.��#��m~�k�ʽI	�){*�?@��Eߡ���⨱�ƐchG�tz�����#�M	�a`~��0m.x��$�%��[�����ş�
��h7�ȋ��2��ZA��gg�JrE�@�]�����f\U�K�5z��y��v�-9��O�B��7�x���D��\g֌"�[��|pVJ��8�O*�ͯm%�5�r��`�w����z+�zA�#b��C*���j�+�p��m���}��|�a��vC���V'#_B�9�W_n9� f�M�W�zQ�J��Q~T1�-?9M/q�{$�ڣb[RH��c�/�͹R�K�Aݗ�A��,�HÞ�(ei`� ��}�M��BH�L��
�P�a������$՞��8����i�,��-���~�����