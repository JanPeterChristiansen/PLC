XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\P[ �
Զ��M�Ҡ+GV;����4� ��Aաb��6($p����$8�=�A�+�'�ӛL?��@�w`��B��G�7��z����<���İ�Q�}�D�n�RۊOgL�m�G�P�e��Vɿ̉4��O�`v��vTE����������	E�}�G�*�G��ó�I�sˡ϶�҅U�|^�0��6�=��p謇kFk O����+>���N��Gy�@�`q�c\8����ԇ!�}V'���sj�`��$~����%N���j���53�<�ҝ�np���;>鸇1*赽9O�!J���x�t,*��F����G*Ԇ�3����)�@�?�%|qk�պ���`kSUEX���ΥT+0�|�)$����O^��-�����b� ��ln�������	<2Y?�$5�jr A�����{#�m�K��Y!I?��{�$��}M�r���p���ұW޽L�f��;�L�%K�A�\KsG%»pJ��:�È.8�Q��'�o@��� ~Q꘦����IA#�wt:��+ /� ���:):��@�T���"��s��~@�/JB���<NG�Y5�=dg: �:�m�I�R��vi㭓1F���?�t�v�
�3bx1���]0���C����F!4��{�=y�	��	ϮZ�ӔΗT!����3�K�o)f�)����1�-
�<��5��ggIc��`"�J-*��*)��ʔ�$���p�ϣ�5�w�c��\iQΨ�+9��suT��=�fq[A��!�5���o'�_5XlxVHYEB    fa00    2020��|����%��d�� �S�&�2A��/95V���"7'�����=ɜZOp�`X!=��7HFg��.��g^F���7D~QA�/6���59�yL�j�� 
��&%�6��B��}`$}dz��|3��ؖ����ޤC�+N+�C[�-wܴ�-�]� +[���Hi���/�>w*�Z���]&�f�H��C]�i�JX�	�}f]��X���e�o4�˦�y����	p�{��t`��J�8�X���<ً���|=�AD�=��d7���8���$���Ht���TQ�ST�<g~
�[z�$�Mw_�h,un��.�!�X�>n�A��M6?�۰ܴ�����%͂HTp׏�*��'�b�$�U����J=:?$M0�<��N8
�����>��[4���fZ����	�����H�@��_?_��M��6,�=����d�Ӽ��MR]Qﾭ��G ��ǇW��q��-�^lY�Oe�p�	�W��b,�߃�\��t>t��t�����JϺG~
�ԍ��^#٭Q�!�V�V$�o/:�*I��,�^�����c�)��w�s&s"�m_
�Xy��m��'�Yc���n�|D�˓6�V��Q+M�c3������=�W'D\�����speχ��\��c���@�!<4j�P��#%Y��<�m�uzh�M�7��s[ߌ{������ѱ��<㬟�'�[޼;�݃)I��_��I0�����*�wT��Q�`}���T/��2��f��iNM�H~r��":�-���+����<6�,.���r��#�(6k
Xˇ�q�lJ$�0`i��^��e~ �a(����!�<�dE5^�.o�1K�(W_L��ꐅn}�����0�gq˗P�	�t87o���Vtǐ��G��'~ ��~zk��🊝�|�u��S�'���?95$��E92�woҬ����C�ѫ?�&��{�
H��Q,���1Bj�Dz��JKZ��'�H�D�u�����>W������j�Z�&H��ؙ��@qú��mr��*]� 0�i����%֢��y7�)�'�Ā�[u��z+��F����($�~{SoL'���N960�~���ב�A҈�_���������pG�ZN�\�v��T��8Y���,��bDL�@��׫z�Qq��=R����7��_Mx����p�c&�N>w�8hA��>E�' S��,��z�>��2}Ȣ�|v8H�\߬����Q�̅	� ���6j{f�.w<��L��+�<2(QO��s]ʺ3~�o�G��VZ��S`+O?���.����本"p���K��
R��qdm����@%�~1���:�e�u,�;�pP�s�8��T�T&$�] ,�&>Q���@L�\=�j��X%4kMԽ���+D�~���j��f��-�nk5�F���	�Dߜ!n��o}��u)C���'�ݢ�6T�D���*�M����Ŵ�r:�,`HE�pw�,�'A����"%�\L�(�ݣɬ���nb�- ��w��ƦR;aL���"�#.l��q�����tm����-a�BbU'�Ѵ?܋`�'�g�Q��M�`�����>Y�"1��F�}u�ʴ��z��B����'yD! "d��3��g��b�}'�w"k$Dd���Hoj�Aq.7X�+D����n��S
�y��"�{��xS�ԫ>ن)7�w�JFj�J�5��>7���H���O1/7�������ʉ����/K��;ϵ�<=�Ѓ
Y$)>G�2��������yk�:	���u���e���W$t�!G�����}'���^��R�Oi�sC���w@�����xHB�Q��c�b�fh����uȹ��8:T��8I��}í�	������G7�|k6��q�_R����9�,7U��E#�+*�8�1�ʒV�z0#�d�k��mh���M�	\�kB4�T��nW�����}b��`aH�U�����4��5<</�Sk"�w[}
�ED�D���,_�L?Rg�˷7c�X��8]~�
�� OG}_5.��;#�k�����o�K����\e�޺&���q7��J�b]�.i�6M����+�-�����1�+N��4��A^����H��q�d�L)zI>�����j��}Juup�4i����?u�FK�w��/Y˴���T���8PFa�;B͟�K�2�NB<�~޵	w�s���J�s|�)��[�JW����ʣ��=me�AM�-p��a��zc��&o�?�9�Q�=C��W%�c�y���J��� UTrl)���CPs�ɧ�Qr8�lu�$�M�ZEX;���`:EG!�6�.��Rȷ�:܋�I4�_�����
�9�Lh�W>�2 PCsaq��9��u|�ZN����=S#O)�l#�K��<��KW�����b��}�G���Pj�s��=d�5��N5�z�B���i����O�[��#1�|�Vh�IT�$S1#a��H@�e�$
��=��>A�A9R���u�����뷘:<Z�*@���/C�?l�5��o���T�����ʬ�x�բ�?Q�O����8Qt
�k7zF��_��kX}��׫7@�=\���$c�?�!2��"�̛�NJ�N�L�0�����ffŨ��	���7��*�_��|Qp�S{I�#�i�]��Dh��Ec��+����z	.�-�H��Z����HHN�H�Ƙ;~0-���b��c�V{��}��t�<�Mh-
@�y��h[��ް�B������o1�_1��_XA���y���f�]� ;�a#1D����k��F���ݤ,��hLpb�&���KV�Mi8�o=�#6�ʇ��6�O�l����+P����+�����3 uH���E����=��0�$��i�T_��Ve��k� ,���e��ւ�gD�v��'�|�<����R9i���\\���C�po��$�+��G�ptb�G�y��1�{�oU�EJx���e Gʭ����N<>K�H�#�p�Ҵ�r$f��]uo�8�i��$���+����g���.0�ɁR��Ob����r�:�\�u�ަ�F����R�as�6���'A�n!7Α���v:P{Ľ[E;Hy��@ �A
��'�#�bS�J*fsk�^};����$��9�:�Z���o���wJ�S�[;��;���r�Hh�ʲ���d��La�yE+'#rT{J�X�A==LI�Z[���l�+����s��|�e]� 6�4	)�?���zI��D'�0	�8�=��Ξ�����:��h�Om��m̑SF�G_�;Fge�	����ld8ŭ_�HA���U�O�3�"�v���q��Y?rRc�5��v�n����w�}�@{h��i0$���Gah�pZ�~oM����7��(>�[п��sh�0꒫e/��6�iN�@l�ѷ��|;-%���v��_f q��B�>=�w����w �]� �h�eU����$�E��&���m4_��5pD�����ǃH�Qyz𲼌�g��\20�!/v����T�9*�,��37�~<&�r��%
��cj;��:|����c��j͇8\��4{�x�#ٰ �y�^�v녟)��]��ɮ �K�%����:��B%���9�i��`���h�����zɤ2:/o��qn�!\�v�ejK�`
)�����u8�L�$���'v��Z�d���ת{��D�q#���4\���#B�!��0O���@F/�#�I�]$� a��P���ԘY��_�<��9�+ٿI�*����kAև�H! ��� �����`G,�N!m��Ƕm�;1 ��Z��Iʅ!O��h�p��
g�.l�r3�w���eN�
[;a��iͨ��O�a�F�(��5���):O�h95R����Aշ��<1��oɇ/�Wt@k�lPf�@�=������o��]��1&� ]�*[�l��u�e���&�1�=Z�r�4;mN֒�CYv�1	�2���n���*�?�h�\�[k��P!��R�(���V�c��Kv��H�#�"$��l�H�I�I��§@XCٸ�m�?$��}��C(�YF�?�`���W|'��خҐ�	�!���H���mU����q_u$>�B!8�����^�)��DaP�pJ>\])��D-i0��pRa±�����`N�;��`;Y�4Vނ�=j���:�6�qmM<0��U��G�ԛt[r���	,=��7��H�{4o��[R(N�Q=��e�ݽHVՋ��4�{��t�E1;"�}�O�r[�jz\{U��zz�c(��"�M��q���:�`�㱧Fu"�";`,)Z�W$3�t�wv,%�I��M�5|�|���30�9/�Q���C��yL'�AF���S�H�|0r�(����p�<t�j��T1�S�I���]����N��k[���M;V�2����y�\f�>5�g�A�긥�g~���c�3�3Z�8�
���{�x�$�\1^ϫ���JI��S����ʝ?0d�|#J�tȽB�Dr��e�[�M�Hw�� I����,+����B�f�Ph�֏P�W݄���N�fe�@Gd6�| �V,�`S��"�{��q���_�f=BʮC����M�7d�FE޵*�wH��o�sf����P���+`3J������zGJs,�Zi��V򒼎����h�3qAd`9G�H��'����(}�X"�u1M�/W�ʤ:Mb5�;��,�񡿯/����aR&)ߎQs���ɷ��h[Q�2U�/0�o2u�����@��l��_�/���Qq�O�{�ަ��C����o��rz��c��,R��,�#p�t,ޤL��rC��
"p>��}����{R�6�O��j��+�+�	<.�'ys�&��
{7=rǡx��ǧe[m�e�v;n��N��3W�exD(��`�5ݯ��qԍ�+/�c�����;��~�QN~�Ws�r��BBv�/YH	%�G�<���\L�8!�s������V����E�*`W �k��U{n���W�:*���GCp��5@ȸ�͈{AF���4j��z�h���n����W�&�ap|t�%㞼j�����@ʑ+j6qn��zmr��	ظgU������
Y�w�$���������S�-��alµGJ���rS���$X:p-[�H�H�k�����l�K�<&�a� 90�3����V�D׭1�b��fi T�e=�ߘ�;���[5��_yL�8	��p�q�c�t�#�8m5Y7d�V5�Bt�g,*�lH��Z�h��{5`���v�0<�[�X�UTϊ���I'�d^��3d���넟Fet�[�8\�su�)j��'����[�ۚ[���@j��ɳ��M�����}2��C
,�}jH�N�s���'oQ�d}5�j�-ωqϪqu���6'���ʻ	����Ki�� �5o@ż��R�/�ܚ^���X>|g(t8�ͺ7�MnT3����b]蛳F�Ɨ��?l[����`�8�W5 ���Q�B2�hNf��7c��r�Q��
5��ѫtXw�����23/�v��� �W�ZM�,!��i�`c]�+�܀��G�P]�;���<��2:�D;{Km�M�Ύ��ʂ�X��8z����ٞS6������ӌH�JbH�)�Ot�kd$a4Y�.�P���;W\��Y F��cd9��&�ɭ��j�=�@Qz��ڣc׎;��2z`��ɤwS}��M$,9̓��͇�?�j�ƒl��z��K��m��88qD�`��vy�y]���z�$sqC��d���Ou�22�R^#w��dym��Vh��:�-����_J>]�L:_abB����9Î-[紶s R��'�w����KU^���X�IXS�5�&j�����x2�\����&gqk�sM�S�s�NZ��!�cN��#�L��
���H��B`kb�5�����g{+T��ؑٻ��HA�$`�����%��`g3"��-��1���:݈��V�؝�w  Y(�ܵY� MG>g��%NK�P�89�~�D7f6Y�c�O6xY��6 ͹�`��C���#���rl����bh_��0]+�]]�� �y	JjL����@���D�Ӥ4�>�:������*	v��L�P��a��ghq�Ct���8춈r�)�;S�!�?ｐ��挜�)Z'T.�Iu�G>(�t�_�Z��3��3�(q7�j,�E˨��!t9��*�Yd���W^��|sМ��R(��|����D$n8�w�`�Oh��9q��I����\��M���|ѷӻ�W�ўh�����>��4��fp�'��.������/��?����fQ1C�n|��?���D1o|�>h&MZ�A���~���np�-F��.Z ���$�S�p!��
[�W�#���W���"
�Ss	BΙ:S�^��xH{LG��'\����{G��ŭQ�C�%�R�+H�x�i�*|qkv����y^��^Zu��/�C�Z��E�{kȬy�x�>�70N���ʬ>�12���G���d�g���h�O5nŔ�u��cQ�g����3�~��w;����}�1�3ˋ�v��葇��n|�uy�9T�U�~��~;��Y����P���K|^+o�
{�K,�����e��T�GJ��G�JT����#9�`�:�^��S]UIT�`��R�C+����<i_��m�z)�����V��Cq�lF�F�s���ӈ����5���?;�\�*Y�c�8=���m<�v��#<�?#3��h��P�Z%4m*ۥ�L�>ˍ=���z���uFfیX"���ٵq}=]��p�=����|h������P#�t�.���~���4�r(���i��ER�R���["����/����	��		w���:�g�BL��� R�#��+��¨k�4�(���=[ǒ*��m9>��B)���/а��;��YR���8��� �Z��0��5L��(@X�=���S`?�U�ʩu�+Ù��VH��k{c��8Q}|ŮX���=��8i�
5������L�Bľ �a�4�� ���������Z�'^�{�i����kgy偼Q�,�y�o�9~#�ۮI:=�q�_����&�ݙc���o�|�X�m&�t�o>�xt;b2��O5�'�6����"d�Z_�����%��K�ԛd`�AxD�,��@ԺY�b��$5%���C�áTU& 9��h3����5�-P���@q�R>��Ֆq���\��"V���
V��z ҡ�7@n��$j)�Xc"�;o����>��h^De��u�j֮ i�6��Ւ7�V�^��ec�U���i�~�@����E�ڀ!0�?��s�o�O$8�=�;��C�X[AG��!_������<f��6k�4[���<=MP�I�J��>l��$8��I3O��j�[
o�/�`��/J��[��R����d��%�J��k�<4J�ϐ
V��!��S����o���+�}6��1��:�l��
�s��J���v��1������gi�A�32)�����eXep�F�&)�;�N���I�~����8�;��J@[�Y��a�����W<[�.wNd�J�6��D�������j����[����3�p�,�dk��T2(���2Q��e->Ȥ�#�8T�o3�ʜ����ʍvy���0�|�Oy��}t��e�_����P,"Bi���_�HNy��W�N�K1(t��k��(��2|
�����z-���_R54��
�u� ���,��*�>beH�ʑ������l܇ �a�Xx}=	%;�ߕ��[�̏z���j�~z����� �J{�r��Jd4����}�uF��:m4 A��¾�g��q�#��
�ǽ�I�HT3��e�(��dfy?<��D����gD��ڍ���*i�%pRT�{z��`H�g�2���� ʇ�a�c�$w��G�c�AS�ٹ	0BYh���"
��*�qɦ�0�b�X����������t:�ڡ����ǋ �0؝o�"D�l��{�b&�[�^V�0�,�~㥥�9�#�9��<z�P�U�I�iݴ�Wp�N{�"�Rm��4L��1G�'|,�t�c%�D�|<{�|�m�7����"��3Z�z)��EL��:�2��	~�VQes�$/;�ΕXlxVHYEB    cb82    12b0�3��o�1�>�S��:��絗7�ȏ5ե\>>��'���Ȩ�+Y�"�,�>p!�;���W/57��i*����`\�26�n �~8��sso�ǫ����S���j\t~��6��p}�J��X���*���b�F��6��,�z"]�C�L�_$3�v���=�)*�GeѸ�RM���z�/��x��PDqv��y����ׯ|�����W�b8�u��G�#A�/݁�>j2ڵ�����_�tŮ��s�a�a����!�k�w��,<7o���B�N_�0�/�U�&@"'urN{�X�J5HpmO�ilG�'�P�i�2����_�sH��B!܍fi��g������G���e�!�7�E�Y�M���v�)%�w t������ޑ�@���E�'R�grR�����=���"W�U
!�i��w�W�V�	������҂���<��Z�cz溮���i�^�]a˨�CE[�9=rgZN=����H0�3zuN����2Veۈj�AW[�Ob�2 ��&i��$��q�ZtD�d��~��;Mhܣ\���M��a칤��ږ	 $��
G]��لf�)�+�n7�C��F�4����Yɼ��}�X�_��r+�t���_3_ze�Hn�U5A����Sľ�O�b,\��Ά�[�AE  �l�3[�r�wS�.���&�ޠmn��'���	6��0l��F�I�܂��FaT�ζ��ş�T~�?R�?��v�M�}Ò���O7�3�^U_����~-�d@h2���bB���g���"90�.�#�lo�1$�Bʞ����_h �=0K����'��3p�j������o���f9Ci��0{�g ��N:�.̚�m�E����M��Ĩ��gc����[!w�o�\C21~�d\��%Q�!̜RA��WA�c*�!� �R�*�����s
�{Q��d֜n=��-t���q2�����~����ӌ�m騠Y��dCk���-s�K��q�e<�K�tӯ�D�W�׷Մuˀq��얌�����VP�Aǵ2�C�ƞ�����	��>��K^կB߉�}��aLy�m��A=^���/�3��X�#b��C�6����F\[�'}��-MX�~�w|Y���`ĸLp��nj`]Z"t�pٵ��K�כ��P˝�/�����q��{q���9m{�	�a���Ub�������C�Ĕ���
E�R��N0]}��t��t P#�@Y��j3'Փ_�<����D�f���?G�b��r�&H���;�?�f��J��LY�om@p
��g�ڑ�Q/��`w��0]�Iϲ��M�7�^$�0F;YZ�В���Vf���j��+����TUyqs���ơs�Lv�<�����Pﾳ�>F�]����-�����g�D@����;Tx{3�>��@qq=v�� rAPv��8?dzA .h,�/��2�Il�g�'W&���E�oo��m�aY����TDmCR�fo�������q\�s����,D�
�l����B�bf.�s����D1n� T����Cl\f9�Ŧ���k��L*��O����E�Da���R�/v�]��nf��Ps�b���mVq�_�'&D��?�G*}�DC}�mPp���C�����B���kN[1HR&vz�g̳[!pU!b����-�	/rM�gSeL7��vȖ\'0��/��H���1־GBGb�����Fħ���nD�ƪ��pj�Q��&I;./�෤Ap��5 B��{���
d:?���z*��Ca��	%��dP�qV����*�y���qZ؄av,kO�q~�>4�z|+zҩk�*�Exb��6K��#d��y�ǙȒ�v��9:
o�b!ɨP0޴LQ�9���!5SP4��g��'dRbY���16F޷��@}B.'F��V�)���	��f����t����}�r�?ya� O:�P���MB1׾M�A-�]0���C���"X��������5>�f��1a[���iU�+yH��|N3�G�����H�}���]�%�CZ񚴄�P\�~���=O�
����#4��+�D78i���r~�^re*v��CV�/"���}F�� ndW�j\6+����~ᙊ}�+�|��0��>%|�����I��a��o��o��ej�>hx�
�&���m�/L���U�T�͆h#B�)4E����kɆ�~ ����`=���~[Z�_86� ��/0��{Yp��h����o��x�'\p��E`�T�2�L�^e���n~Py�l��?�K���n��7���Db`�x[�#��HR,� Xs�	�^��@
���	�K�²��`�U%Y}�f3<�
��&���$(�q�z5,j����h�w��E�	�?�������WT��;Е8�q"
t'1���dB���AnD�|��ʦm5��W�O�ቬ	3�j�������~�J�T.��R�5�ә�U��P�c~��H@��Ys��BU�`��Q��cО~~�K4�c��(Q�� 5�TU�Վ8{o�p�.{06�o��(�Nлe�}�s�[�y�շ?��+|8A�
Ǫ��c=�)0�Mҝ�䃌��ޒ���Zn!$sF����:Z�T)��E��r[��A��a/`Q�FA4U=@ɜ~�~ �,���yS��^6�G�-��`�8���u���`��up4K����7�%���rp%�](b,�Z�D�p��x��k"�; �0��Ϋ[O�W�����ж�@��`?��/��	u�L�y�9�ﭻ̫��r=�$$���.X��iz�t׿�z�x;�w`�n���'=���$�5��D�{o�BE�'�@%��|!�*"9LϮY;eќ�<'B\�2��ʊ5�Fft�'Qbio,���U�Bpn]�n�:���Y#�*�}DV�(��#�k�@�t�u�χSJ"��M
tA�*gz���0�|V&�������=�1(ӡ�
"��W�	0��f�����=�{��>!i$_�~����]1�� �?�A�����M��E �e8�j���E���B�w%ec��^?��{��n�n���_��k��/�� ��0z���\�WUl�x���L�z��4���V9�7�Ϙl���ΌL6���<�:xB��iH�̔��%�����L:�+rȆH�6dy�9�oqJ��\�V�1< �)}���f�ϓ�eo���nH��m-b³fs��ڱv���R9_���h[�ۣ~[Rqe�o'�-��A�XTVG�ɷ'B��*�	�N�ӕ��"q*텣�U��U�V��N��A&°ԉ�h��)cqOWͤ��t���#*���~�\�4Ӕe����4x���e��\ܙ,:���Wf�i��+\�{b�QE����L�~�ɘ7������{��d�ԕS��~e�1%fYMAPf�9�T�ݢ�&/�[���<�Ԁ\h�R+, @?��P�C/��A��~_<֋����)u`�~�m-�g�ۧ�.��SP�rp.�&Kp8����-�(pji��Χr�C?�wD[ �e�g_/��}ٲ���_�J�FL�h�ޤz��P����R�f'�d��HO��ap��I��$P EW4�?�����L�F8���-i.���� ��[���<*����ÿ�[j}��{0H{�{�L�1}���3-�E��.wk!�䍼���p����١��]} S/�&!�l�ށְ��}��l�tG7��I��%�s�%���tw:G���y(�<�a�&.�y�:ZU踛�gܢԶ�gv����g@�iBgGvR0��b �X�*3���Q�N������U�DUB����Ѹv-k���7$)�\���g����K�Z>�)��������Zv��_?��aS^���>�/�J9\�_#���Jh�<�����#�)��Pڷ��K��eU��77�(���(�xM�ȼV��;�֛~���Yt�T��2C��K�QB�q�y�m>e�m�����fΩ�xX�z�j`��<��#!�uJ��� �>��N�Ed�j�ع��`"��J�,c�l��*cv㘥�=�S������x�(�5���D�P�?���b���>x9.�=�����\[�*���n], �S��V*g� 2�@�|e�3h��d�ޯ���.p`?�d*�{c��OeAζ
�k+�����0�ǖ'ա����?���X�drCZ��<������Kl�s2 ��XJ�/�����t���.�{�)*�B�Sh�[eu��y��$������n��gca �*�l��F����g�ڱ^�r����'�R�hM�ZMhn&�Yt��={��d�_y(2=��*�M�%!\��t3���y��}�c�ĉ{���S�ܿ�����2�iZ6�
�5'ÍAd�N�Dj	Q�o�%�ˎG����JV9��*��~�J#fO�h�b�g�[aH��������?��~���Bl���b#��a_��~'c!����!��t��T��9��ai!t<琪������%����D���*���˖	O��3竖�K�,�h˼1ٶ�f"�\��;�,����\�7�Ց�`a���8D�Ty�Yn74���|��T����=>Ƈ��X�
hQ�ntw�P�.V�#B�#c����ɌEXgq�`�|_���f�\�d���Ng��D*	��?����25k*�.Nh�e�UGiC����4�wh�eR��(�--�V�ᤪ��k�^+���9�.���������JX�Z|��F1��Eຸ3l�