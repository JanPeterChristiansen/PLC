XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ax#�\5�f.}�uy��x�L�!2�;��>0�g�=Wx�0�m����<x._6Oj���1A�#;���,LM�tm���&R����Ƈ'��,ܙ#e���I@�?��K��3S�)���`U�U�+�'�O-x[�
�;����� �T�
�wcp��1j�-�� �����x_z��΄G�!�����d}N����c^��{^��웮�`W�� ��5�@&I��������%���+�
�C��T	Bލ[�4fD����dy��T"��\�-���6i����_�q҂Ֆ�#��,V-E�:����U(:�l.�	yx�o�׸��Т	�z��oĚ0B�r��*-���D����<����VI� �=c�y�Dy<Pú�J�#E.�Z�$j�=Z�w�D_��0,�����56�<�t΋1Ѱk�:Mć�KC�{���9<���Tq�
��0�V宭��@���ߜ���:S�]Oq�u�=�x*���WK�ӵA0��z�Z�/	M:5�O#��.���Ғ��¸(�M�1�f��PS�9�1}Jajtw��p������*	��~�˳Q�Ҥ�c����{4xE8�g���lDq�5�K��h�tK�f�W��ș�����4@f^%��rw�^D����hG��T���Tӥ�-"����5���A|�Z&�����K+:�&z=5rF�'��e�*�{à�����E��%B�ADqD ���iW���F���XlxVHYEB    c3e8    1d20@��!Jr/���o�%���za����$�u|]��G�C"e�����p���<J,'�7=<�^9��.S	k+���_�J6�<�R8��� �Q�$Ǎõ�6��c�,^V$�T��8
��?I��3ql�n�^$:�������&�]��h��\
J�5���7}z���a[�J�[Vo�l�n(�]^1i�5$�fP�j����΅�o��jO(�:^g���F7L}��*'Dؖ���/K+�˳�H�Q
�Ij泉�ݧc٘�p��;40q"���g$p:�M+�m*��t?
����O�L��
s`ZD��3 ����<��ʠhEi�ĤF���;���s�������B숳���.Ăs���_@��xܢ������0�{T�:�*�]
���gs��+kYAj4-!z��#��_�m��v�����)|k�~�������?�(`*yd���1xd����K�|W�u^MfĤ+���U���4��S��{��{$S�S�:ƀI%��!ÛT2��<l��kȺ|FJ�t_'�����Sp��������%�ad[�T!1,�'��.��JަH�20�L��{���/�2~y�m3�nʉ���OR��3�*�K�sQ�SD5�Kz�z{������^x�kɔ�CB�]"���cK�.V2b��}qf5[�4k ���5���oweF_�2;5�����C$:z0�W���"ퟓc��p�&���!�|��@ �����p�u���S����J��[u?.��"8@˥2܎��-Z�ۗ����#�$o��d�d�QcY˒�zm#��U���r9�w�E���:��ɪz�������b ��:��EI��;	�s���wI���#�ӎ@L���NU�3'��`�A��p ̝�xT(��/~X��b���>b�z�(�@�1�nt��V\+�dr8#����0��3w__]�j�N�.��e�	��s�;��x�s*�ʿ�F��
G�U������E���@Xn�+��$f&���xa!�h��o�U,�o�]�M���A�>�� ����i�5��Б�9��V`�Ŝ�Ѫ�wM�dr������M�D�"/ޅ�}Жqnu�P~j�g�U)����	�:bF�@ND�X�P��Ԝ��)�gE�l��@?H?E�J��,�#A�bY�����+����o<��MJC~`����3	YV|�ȍ��t	`���*��M<�=�GmYl*��Ӥ��d��a��	J�-$���h�kܻts�[!�T��l�$�� K�	�s�$�5kN��;w)��2��;���[��:���5MME�����ʌg�kcb��R����ܐYqk�� �hr4�G�-n������ׁ[�,l���m��2�63�N��-�u�u �ɟ�����۞׹]3���bG��-B����=���l��J��G�x�O�VVPtH�D�ٸa"��ϐ��'fJ���>�l*�xG;V���p��$@�]����L[O���isp۵�0b ��[�r�WO~`^���ً�1��
9ڥdp,��\R�g@��;U��QvE1��odDʐ�޾����?����p���&�(���*Yp`��ѷ�qwׂ�4u�����&|���꣉�g�J�P��ѻ�)�"M��kR%���@"j��Ѡ�QS��P�,����N-?ӎ���+&�?�kA�^�,���n,Z�݉�V�/=�=�ɷa�?,@���t-M��_j��_-��ZPм�Uĭ��@%mN��O	D���yT���~�T+�2%�u�`ʜ�G���v���j:���$[W�$L���9#G��T��ZFEj(\*�V�	����b�JfDO����$&Y�����b�R�ɦ�7��l%Ҏ��4�T֑���B2�H �-,+H*�=x�sj3��_u�T~3'����?�=:2�k�0�G�S뗘W���W�7/gc ����X�$�ZnJH�X!���`me�	d6J���$O5hi��K���� �/��y/�@֯���qΌLܵ��Wu=�X���m����}(�E�*Ð,�U�3K���m������5�X���M����J����o�h:,arۖ����]uľ(���?d��8��<-�[�����n+���؟��Ҏ�/XF��7�����cE��^���zl5�K�d���n�8�my��7f�d�8n�H�m�?i��(�r|�]�[���tC����q�c�s��e,�EI�Y�j.�Xл@ԋ��:Y��7�C���`R�6KQ�DTd��7c�nOV�� 1F���GڎF���?�o��jnx,9��|���~�V/����a84I�&�iB�le�>���b-܏ȱ1d��C>�(Oާ�N/9����T�M}2���7s����R��4I.��VM������B�n��UgJ�<d����E����sgfwY
e�|�xЌh����o�w<�C�Z>�X:\2�k�D�Jާ��N�;�����UK7����&G��yLD���Gz�]��Y�љfp�<w�ޑ���;�M��vt�j��(+BQ(s��&��f�b�q����l*�G�g���YP�:]�����|���p���R�$ ����B��Y���f�������e�9uW
R=���=-���+l���R�4��Gf@gJ��ܙ�P%E��y1��4���#��5 ��dP��~���ׯ��C����ӖUMzLƟA�����f�� �6�����)xO|�fՎ'JPo�8l��ܹ��ǤrD��It��7q/<��)���}�v,I~ܿ�gX�OJ����ґ7G�!����7M�B;�׷/�2��-�ĳ���gHա�4T��	[zo��-◡W3�	`���Q���WtY�A�>�ݟ��&"$o�-�nf�a��9g�j&��US �^��|a,�DON�ټ�?��3�?TC� ���X*r�Ә e���g��h��D�K/f�>��$+��N�Н�%�d��Ѡ��;��ՃَR�z�8-"��[ۜl<Vhij�Ĳ�o��t]T�#���0>4��rg��(\�ѯ��#�ʫJ�Z���-�(��S����.���*����hԪ�moC����K����p�0^��� ����e¬n~�<�{"����QG�=��� �gn&W&��<nA�^�jE��Q\܎�XϒF�T���	��9�k��R)�f���q��Vu���'0�b����v`���]Y��v���%
���Dï��g�y�7K���M xyt�w�l�[I����K��6�ϯ�:�M{�	�	�.�F�vET������O�|�/�t��w�.mϗ�0�*&�����q���"_zs�`qY��e&���9���n��L�D�G�� ���?C?^� ��-�,^�U�o_�[/�[X��Bt�k-R��e�J�֙%]E�]� ������{��0���\�.Y9����vv���2��H�ݥy�[vI[��t�dn/<�t��u:�tEH�C�R&�%s;����Rb�1�������j�4���:�|�����f���\�:�m9m�a9xK̢�tG�m����j�y6�i��hH����}�4p+�~P��I�^�C��i�&mM�cej�<si5)!�"c�,F���ɒd��Y���T9z�.�1J/�k��B˻h��B��mEH�[�sq��;�{�W��V%���d����YO��!���D�"�����s��D���a"+`�I�;�
�X�1@<R��Ms��݇2�`4R7S��U]]Ü���H�:ziu�ȼ(���E�HD��w�8Q�	/�O�jlW�Z��y����كhwTW��塻=^����Ͷ$k<R�2����\�h�r<4�d I���.���9�jq��aX<�)�⃘`�v*B��1R��J�E�Vᔯc����x�#ݙ|����5�j�N�:���d6��'�56`@�����?�>���Zվ�%~�9�׸�y��C$7e�#�>hc����=�w��R�g��ތ����	�^ƶ|\U��a��h���:�_���{��Ƀ^Ɓ�ncw/��v����哞F��+�GG:٢:�k��C ��'Z�&g(��/���oKn\m[�y<�V�L����e������!��QV)
�Q0p��ԔK<ځ0ذ�^n:�s$F60�C;���Y:Is2��Їg�XI�2I�힖�9�S��r6Y-O���[���j��U���?"��"m:=e��!������- <�h��7�HȚע��<AJ����C�O���!��^
��)a��l--��mg4�`9f�ZtN�y!`���Kv\J�����,�!(�4�J�kܪ�I��YZԘ�*�Р�1��iv�*�J�H��N.^��ȯHL�<h��A�����wq*'8E�W9R�-�m%�ĨK��u�X��<C�b�m��^����T&����W�T�}��jj����0H{�����Z�]��-�}�zu��3����j�Q�Up*l�Z�K(��l��oZǝ�=�[�}��r���,8K�!7��HKuӠ��`���TC�A<��3�#�0���95�JI��+�Ш�<�p�m�ŹT ����k%zZ,�.�R��}�t���Q�q�azQ'�d�IxJy��<-��P(eñ��� �d�%��cJWѣ� UG�cX6A�*kH>^`�Q��Iұ�p�m|�ǈ]9�W7��6��0���IWp��_Ϧ�إN⧎D?.�y�x!�Rw��ϴn�a䷳��:����~�ޡ|8> BK&hR)��+���#�eQ���8z+{�B����hs�����Ō�T/��y�� � tW��l���{�d�t+
Sa��<����r�7aO�h��Ё19j�?�N�H�6]�C�d�$�}�8�I��&s�a�M-w�f��J�0�J$]_I�K�^�&x���JG�`���?��y>δ$FQݒF�k"xX��}��٤�9k�4�����<�~$���:jI������.nb/�����N?�
��:%-!�n�;��mhs+��j�BV!�Z��V-x��慃��b�e[����c�;��k�D$�v"/���xD7'���[��i�~��ｆcYH�̃@�<4���3U�l�~�?��u�r��������!�Z�-�	���:|��}Z�~�p}�|u#��fՋ�t����#م�E�#q��� �OMDUo�k��?آ��)G�ow����0 J�����Y�_��I�l�؆:�3�U�)Lk�lu� ]��<u"�=G�V�ѐv���%�{�f܏�"����x��c�L��5'$���<�l-�A˥7j4k�D?�َ�xYM��Z�&�'��w�Q2�O��g�Vӥ��>5�-)�p`A`�����+Z;��lc^�V
7�m�=�����[�ٲ|Y�2���G
:Ҷ��N��� �k,n{8ٲ�4����LQ�m;��_RV7���]�����3J�⃦�0fm��i,�%�g0{�wU�$,y�M����Q�z��I�8�~����W7��=J�;�6w��6�D�$�xT./F��@�'�%�G~���E������
No��gK�l���V����LF�իYл��l�{gw�z�Z7�n.ʮ��E��s�jd��\׹�yg���T��zu�Dz	�X��C��.u$�T"SG���i��xǎ������_pZ��]�7٨^����|��ܓ������p5�#
PNp��$u�~�{R���͆r��ݢW������lx�j�����.hޖ��i� ��(ّ�"�Њ���n/��V����Y�\���r"��q��a5�bȶ|m�l6߁�$���9��R
k���i�rZ�Pm�T�6�&��&�K��cw��3���+������yXP��~����L��RF{XLII�,�X&Pv�c+�~<S^K�,��ّV<�d�v���e�6n,��a/t�[����&����_;,g���K�+���J�itLS�*6$���E�_�r�U/;_gڧ�l|/�oE&�w� �����A�~�9��w�ZӀ���@r����d�S~Uz"�t-=����Sb"?�j����ɞ�w��9t�웥6�h@c�<7��"o��;��p�m
�ꋯS�I�a�`����63�#X71b%�μ�{RO�}��8��9�c���$I�c����=7nf��33,v��p�2衩����ݑ��B�� t
�B0����/n؛�<��.�8l��|$y��/< �ʝ嚲�;4y��q�!Wcݻ�Ъ�+{��tN��F���K�kW��kVGmP�B2.�t���Ӄ�Q���Dd�#ú�)z�i؞ne�?����즦Z�^��rk���kK���V_͠!u�fK|s�m�j��'��~QǗ�>e�(����o�*��%R�y[� @Ò���`���@��K�ݡ��EG�#��d����lU��ڇn���|��U��f�p����L��&�S�A�n�OI²�{�����4����g��r������"��Dr�Z�4����vl'wn!�91���<6P9��Sѐ>]]�J	��H��BbE7����~7��*��}�T�C���λD
����3�1،Vz�Fn����x�$�0=�����S���j
\��L��+��� �; ��0�{�����܈���܀����u+��I��H.��kK�b*�ѫ�?������c�"d" ��R�<_(�5�
��_�-���@M
5������(�1�����M�^07����u'�ediBҢ���-ؿ��\O��u4��a�m�:c*H.u�.���,|���e`$�}�{���i��^ƺ
�k(E����_:��T�!�)�~FL�f�w(H�\����:��ײ�M�����7�
����M��\�4VE��v�\é0zMrc#�4J���ߋ�9G��KU��L�NMq�A�.�$)�ka�kL&������N%\��U��H�$��O}*������$�F1�w���#ߚ��ee���u5v��!n>���l�fm�DO�"�H^���Y4oӴ�����f�*��<��2q�l7�#P��-B��"k	�;V����"�y��6YAT������;@�Z��{i��9֭)�*e��E��(�Z�1���}���ب�g����.���k�&��� �|Ҵ��-4e	͝���Woh�����{j^"+j��L��Dɤ"a���t	~*��Q?R	<�=�|����˾t�,�{"���g�+��Lc|>������@�IR9a%e�ұx����_�-�Lk��f�����ކ��O6i=\�����a�Q!��Ō,��w�͑J4
���>�W�tK��(�>3��@���