XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��n�\\�=kKRn���M���R�M<��!\��%���K/ԫ�h�_��2J���
 �<�d ��^qU��x�K
0��dI������ah���Ot�\���uyG%�I�K`Cd!m��
+�[��$o�!#�r�"�aձ;��ŋ�W9�P��2�ۖK����P1X�?F�J��r��D4��ֽ��K5�C���enr������h���j����������@��toC������F�)�`��>Y\�?��&=�xo,�x�.⓾c���^Jm2g����E��*sȌ��|g�._[���&�|C!n5�8����fe�@�t�*}K|Br?�i�&{�q�'Y+�y�h�����������2�Y��CzSSW�[�5�п��Q��:W�Α��^�a���#�ʲE�'In�k�=��C\��=���{���"�X�*0� �w�6̛�ZWT�V�����6"&�$rFV���ʣ_��m%���V��f��f��NAU�J�����?>z��j٘:K�0D����-��X�!3�,.��5�bk�v��8�4;˻,Mj�X�R��~�2$m`��=���o����Mhe35O�ZS��OS/:���<�hs�T�/F�,�Pˬ��f���vJ�J܎�Ш�n��=ҟ����d��ж#T�=QՍ��}_�w��.
'Ŧ?�>��z���}��Z�,���y���ML�i��@�� H��� +�2S1����a�|Xoe_m	��.�-I��?�V�p�XlxVHYEB    fa00    1f80\��Z1~�=cʧ��`���k��c�� ��pO�� #A]�ZQ��P>'�1l]%��p(G=��[;h���90�}W�
���o�zX�l�Tؽof�8A)��0%��>�^E\���u�-��k�J�)i�c����="�<��=>k�͙j��e�?mP�p�
ЀC"���5\���P���dSq��,�N��Od��!� t6]Ň���=�;X�����*�Wu�����r���В*��nڴ��Y� %�A��%�n��0�"ژC��I�|��iG>���ʹ���&� ���.u��*��aj8y{��Ɍ*F�獞����&r�����.��aOͅ�{&=��d�����˗LaDǟ���pPƊ*e^��鑐�,�z~�C@�+@����{��5�Լ)��V߱� ��q�V��J�5'���`�x�9
z
�&0T�X��J2�?o��F[cx�������a3�Q����	mUV;�	�2-�F�ǧ��!�o�4��s1��O$�yZ�rw��D�@WnG�������E�a�m
m����&g@l9-�:��qH��K���B9r���t�K)vأ��`����4W�@�m��f,vI�\�o�{��=$BI܉�ڟ�����Ƴ�7I��zS��/���Dm���v-H�����7"*�:n��p�2cdG�N)��*��|nH����iƀ��'T�mދ6��.b�E��8��=�:8眥'S[	j���,�k���!HR���/�hC-[�1���<;Ʈ�!��5�����lT7w�5��4������&����a��h���"��_��U��˭��i�A����p���^�;���2l�h������`H�W9[�]Kn^��幯����X~�͝��>�E���!�}f�)a�����b�	�n��)�r�ɼ%`<1u��WLe�Z�䮤Kx5�D�6&'�L�R���/5�x�Ҝ��կž�Yo�Y˦�I��M���~49y�K�j]�bH�L/���u�Ǒ��a��}��I�ښ�+���6::g<��h��f�M��L�� ��'|˺M8]��&b����vhO�ӛ���ͨ����v� s�����c~$�XjM)��W�pB ����Wd��4;��@`������0�}�5�R��-���ض�۾I^���{�������読�Ї	��V�V굑�M��.����A�
R[���a]4e���G��A��mF�����f���l�h5����2Nk[N�z�{%�B\�L��b噼�MƐ�������u�A�`�=~Fv��l@=	�,zvJ�r%���4�������O�^�Ȱz���ȑ�66�4��x��CFP���!Ŷҿs��s:�+�*�%k�]GQ�6k��|�Kb��Z� ���7s�m�*Ӷ���64�S�lS�JU=�a[UQc�i���v�q����û�Zǖ���ь������Q#Hk w�{�_��vX�%0Dx�]q�`&�"B0�Y%����-���a3����i" g��ՄT�k��Zf�i �g���U��g�n��<�=�k��a���3)���$w���;��2�Z/�m��`P���K9�w(a�>Zs�[(�qs���d�f�/��A��M��g����q+��$�_��,������6 HG��{;����U=]�����m /����'��I$����@���:���m~�-��L3Ԅ[ZS>�ǉ���[����jƽ7v����!bXAW0�Us�-�ˎGC�aNu�/0�j����.'=f?|5>�E��v�X̔5��0���]����9R�$A[�v���>���Ǿ�h@����ns��,
�+�1	f�b��QQB+^e����/�2�h�my'�S���:.�p�=]�����u�(�qH��l\g�-zT��E��[���)0^ +����G�-|�bϵ�!�"ō\j��ԁ��p�rX�V��3����ƌl-N吿Er����&��p��}bQ�u`���;�We"/�0���^�&� #��ݗ$!M��f�b;u䒯��܄�+,DC	닝�[{).�X��}J��Vf�C.]G�g�H(����+��TO. �8;n"E6H_諒���a�'��ѥr�Ͷu7�5�?Prh�*�$�+�#�1����d��{
Э�i/���$"�V3c���h�?3m��cD�X'�:"2~N:O��T۴�%�[�b<�"�P��m���S $J�zdDh���<��a��%ߏ�x<ɖ΁�ܷ`�fq�y�����F��w�Sx�]��>Ǝ�v�AM �]hΓg����{r�B���M~"F�;���4~���ޢ*�/�W.y%ǈ��9�*c�����ϊ�6�ҳ>PtoF&9��D;�\%����CK#L ]�<���:.�l>�x>Bcl����9αV6����̏k�v(I�c�y_v��}��nP:bc����O�
���K��s!<���9x�"�~蒓�$r�^x���k���V�wm|���XX?��Cr/3c<���Z��P՘س4c��4���✏���W	2"��-�j9�K\�_SD�zX���_Ҋ�Bn�� �Rv�`���R��p����sJj��3I��<3���/��y��s�C����tAt���.la$��J��ח'�ɓZZ�o���҇]禦w*�=P��޼@���.������2�=���mM���S������sN���3��m�R��v�~=�;*����/������;�<��p¸����B��tQ"Xo�Oh3����$f�����B��/��S�����ىeJ:����<�|���I�I��,���D��o'�ד�c(�Vu������ߜ��[o}���f�Y�R�x,����T=y�����=���ϲd��bhP���S)��ζ�LŒ�9�����Ǥ��s;-n\�q�&n�<�Ȕ�'R�M5���( <���n�*��oِhG/[��O�0����à����#Ri�A�e|��J_�z��:�6_��'w�N^��X��`gl�@�����	X�6t�*\)M�#�.EW�L'��I�kY⌲gƀ������8����(&S����7-�ޒ�^�MC%�8��w�|������Eh����|�jET�W
Yb�ݛ ��u�l�|��`u�ʖ�	�W۸��_��'7X��u%%�ɱ;���}_9h��W	H�>�v�T����#���=V3.ş�b���ר�b����	����ݨ��Y쭝ۥk~N��{��}�ځp�P�����7y"��t�SC���ڌl�l:8�Fۑ4�-�3fGlW��Z��
p�(M�jW���4L�� %,`�Z=Է"�=�@����Յ��tU�'u�~�E��D[nK+3oc"�T��`�4��P�^{##+� �c��E�<��.H�J̳�6��?��DO0d�h�� �U#�6��զ��l�4vf�;�"S}$�X�\�b�����C�TA��,L.3�8UJ!V�V�7�.�m.���)'�7d���<m����V��?0eO=�d\�,�u���z�����4tF,�:M�t�at�\�`���]��C�"T�BaUs�7ȥ*C�Y�g�����Z�e5ѿF�+�@��~1������~x����O�e�����o��0�b�a�"��[>�����1EuHm�:�U�4�$���+��Z1�����l��&���N������EuO�3�m� ���#'	�GG��i�i�sr����Ϩd�����:�|����\Q��� �<<�#+Es�5��	��~�~�*��Vo,�?�LtiFD�@��&�İ).�C03`��`JGN�}�t�e�Y����
a��� }��_χ@p�����o��͛�R��Y�<����h�s'&H�6l�+}T�b��}f�:���վ�:��Z�U�fa�co����A;�E_�ίe"��~GYʤ9}I+�
��K�^��C%)C ���I8��f� �M�����s}�Y3�k_-r�<R��'/��n�� ��,!�T��/N�Guy|�)y�-��Z+zQOm��S��!�J���:��V�Ӳ��|z?�q��]�#P�\iL�d$YQa��*�����_��<`��	�:����L
�N!�������BL<l�B�6�
��
^��EI�I+� O*BuE�����&h��w�c��H�M�k�A#n�����:��B ���&�[)���������c&	j�]#�&4�y��NF	Ŧ����W�-�|l���g��kV��d�9��_��h2��7]�3��a�3:N��F��\Ŏ����S7���,U\��ב����f1QNC>�nڂ���<��;/@DH��)��\�O�P�dr������13w��f��Xo��IV~�Ll�I�~��z�
2����EI~�.y�q��:/��E�Z��A���B��G�u�N�0�$�3��@������8��u��!�fG.�Ӝ�Ξ���D�b7����4.0c"�L�u�d�M��Y�0G��1�������γ&t�q�۳id�T����7���U{PC�:;�:�u5'r$��FN~��D���`𾑈�@�8)��\0g_�����ٯ�YEM�LB�`�еڣ���!l.��j�`c>�2���b"os�Z9%���_�w����r�:���'�I�P(�`� X��5~�����FN�Re�n?D�fȃ�޵?R���jJ<��ø��C���!���X��Y�����7E�b���:��1�t��*�λ{�;�1¤��kA����"]��39�}�G�����3�=�=��������5)wU���>.�y'�#d~~��%K����JY�Wz��!Y�?+�?b~,�"ڦ_k)�k�6wk����4�,s:�Ι!����������:9�n Ņ+{���+Z�:*lG�HE��>k���O��BBI�T[�gM�O�R������egT�)����Hu7L�S����
ȷ�q`v΋5Oϟ0(��	#�.�7��&A�f&���s�Q�����6��-)Xk`�Ə����Z�8#����+�u��hoC�'���Zt8v�E,B/:���lH��feRMlWsB�)!�u�ۅ�
��_�8rq&e,��4��$4�����̜�Wj?��������@�	�G)����4`�ݡ��݃C�B���CК� �p٬A� u����,�o��5�l��X0��HLV�ox%�{��E��S�
+-�e-�Mi"��k��ő%��J��x�>�#fT�r�����bd���sD��4a/��������y�'f��WM�,Y��s�?�����,e�бc0\�C�й�髊Ő���.v�z$a�pb�=Z�-+t��F$"�,��M����K�x��bR^��>�X�k�h��%��:*�o��c��8YY�(Wu�y�-�w+�P_�Z	�E��}T϶M�p)}���*��]�6e����7pn?*u�
��QP;��'�ÁWy��*��f���9Ԗ��d�q�Bd�g�̈82���}�N:E�P	nj��^�V���n_��rҘ,�o���:X e�o�bY|4;ol��I��CZ�'(�yWOm��4��.*@.�����a+@2�8������A�Hu����g�?-^��Z����̗`.�o�C�2��p�>�ｫu��[3����V@*�����+�,}������:��U��2I�y��ȑ(��a~�X�ˁϦ5b��T�[�?VȢS�q�#�����P� 4�	&��"��r�W�.Ub&L<V{�*�>�#��`#�H�nD1���&Ӥt+�T���#��)D���ss<J�="5�op�����	��IrZZ.�)�Q"�Ɂ}�{���9 :��!RcsB��gcl�����"�3㵧.����"�e2��!�b�YM��#l�z���
����&��;�0!�T�
���K�=m �s�b�}f�we������1-���V>g�ꉉJ���^k��:֎%G���U`�6��p'vK��g�+�]m,�5PP�กW\���+<qd`w��T�)���y�ڋr�P(�&U�����DJ�o��E��v~�9|k�����}�ҔY0m]Z>��l(��Z9�Q6��U;��W��p���m½�ż2q�]qW��|N����݁��//�9%��+�پI��L
���V����ze�*���>O����ZvS����YL��!��`�B��[�!3L��g��������6iC?�G�4,5�-���!P�F?�z��e���Y������΢���q���Ko14�i�.6;]y��e��^i���m�3�#����+�*�s���L�Y�9F��} �%Šev��A/��g�(M�}�V�5�g6 (���f��ڶ�P��B�ͻ3#a��:�{�2��
���,-�mLk�V�7Po�kϐa�0� �f �zǋu�4��ۉp�G�]-�V��1�%P�U�?yи���Z�/�_m�&(��Gq��]��=���*a���r�g���Y�Ζ"�ID�]X6"
X)Yt%�
��.�m��ٔ���(J�P�bl��jF�%Ņ�����P�΄_G���^��/BGԜ O�t�{��"k��b��gx��>�������vS�*OK����+���~ֆ7�mxi:�3��+A���C5�Oe�깬�f��aX���gl�`�.B���E݂rx%�Ū�{����������.r�޾��X(ƃ����O���x�+��C��WPJ�s���x�a_A	�_���M
i���
�ߙd�`Od�g-7��KE��]�H�1D/|�*<;O����tH5^cư��p�]/��`�?�v�v�]�w�|4�ä��V֋�۹ՙ��3vWҲ��Q$l�؊�tb,h-�7�����V��"�g��	�� �3-چ�����ɷ�I�{~s�Z\ �0L�[�U�xDF�o�F�����{�]l�}q��?7'�Y�O�����S���p�g��!�Iuջ'����������;�ax>��dO���Z�ZD� ۜA�s�,F�׎ҟ)v�rb��nj*Iai?�}Z{���^����mr���k���yh	���E{UDy��jm-�3���HVK_�#�#����i���m�7v����@��������У�:�q�����D�#�X��,�^qa��R��2��0���P�Q˝"W�Ќ(Zn�������c��Ē�*t��C��Źli�!*ě9��d���+��.li��e��ZH��r��h�l�V:�+W#�U����4��NWU�?X�d�n��R�Z�� *cʼ�Vݟb@P	�h����&���\1�.¢�f��^+�����)��z'��T�5����E���rmĿ(����y �M)ߋbƠ>��e�62�9�c��v�L%� N#T;�m�����摠T�(���>AW8 �2+�ȉ��5-�4����B��I*Huj�ߪ��$/�7rF�L�?n!�螉4 7Z���o3�l?:�K�l���Z��$������69qds��{�]RHϮ��ܖ@X�:S���F�v���{��t���O���H����G��*00V��TG>����ے[�f��5�֕2�T ����Y��v��S�U���lӥ����*�s4
�UX�?WU`�
�B�y�������J�mDz��.���������Ag�S݀�,_`�՝QA�랛�#F�,4̹N��V�Z
����ɖn���2>R- u��|��J�,Mh����HPt�Kax)��,��\�C���f�>s�$�/�ߣC��$ �>�B!O��HT��4��kG2��H�F���9��>��]J/'�����#�v@|x�h�(���
tL5��h�XlxVHYEB    fa00    10c0�� �.�x5���)�Њ�2��b)N�l�]�`[ȯ����'���z \ S����뒃x��S�:�Z�/M�}�͛�K��$��Er�\�@�qK0��i9$>�y�2>]V�V
�ާ�?��9z���|v��.%H��\0��� s0�4�عP�ʺݮl}�Y![b*ɐJo��c$�Y�,�1hI���+D8��D&�j����79.��M9����te��o��XAH��(�j���%W��ךxTu���Ixh�Tb�Wr?H�r2c)�-�pXO�cm^ڲ��2�IFx��� `��$��S/�Y�</����,�9�	�1�{=�`e���>%���n0�Xr�{NHK��p��G�����\ �:M�;�;���B�Q�~�v�8_PR��+i>�ab����쫂�F�h	W�$;������֋FvWx	���x��'��c�v6}� �������]�/��Ʉ��[+�a�_�����'�m�>�z�!�S��>�)���xGd�jQ��Ak�/2
�E����Z�KΙ����ߣ{�e�tF*��o�xS�H��p#R�q"�	:�9�˨��S,�+Bb��ێ;K��x&2]Ѹ;%s����3����=�L�:�-Cp6��L�������BU�o�=��v��k �nCW���>�и�� �y����u��^�4VL����Ϙ�����;n_�5�x�N���_������P����g�X*2�no���RY����(!��e��5q�ސ}!�_[��7\���B +�@e��`1���==2�43��\^*'�o���g(� ��k�G�i0R�@�hy
ܻ�?M8�T8ӆ�Tt�&ΥY���mA<�tT����l�M���MO#�V�(�Gy���|Χ��������r!�i>!���P�(lQ/�E��As�u\S?r�G�l禞��Qd�<ѐ�#��'�E��!&�~�G��L���:U�.�������/n5�l�b|�N@�����lfݱ-�E��o�O,�ွu>�<�ܙ��>K �ŧ�V
�"�o$��x���n�d����S>Ǔ�XϮ����7֖5o&ro�n@<��X=�y4�b�L���a�0��,>"��9^�ڧp��~ۯa����b�����5"m���d�]Lf�=���߈�<]��c��N�!�9�����S���7�obAz�X�h�:jJ/��VK���d{3$��>��Ws�v)�pGҭ@���K�����>߷m�_�	.�����cX��wպ;<<�-*�U��:�v�	�����0p�h��W.��2�O�>vp3�O7L��~�ne�������C�鿷��e�����m�r��/�q��j(�+�f��|�i��츑��:b�u�
��E�ح�'�,Q�9�yq6A-�-k(��{ݿD.���B}%'6�Dz����nAȆUr�����v�g1�Y����ԙY�HN�>�Ѩ7�a��Rw�m��R����-��d�;xd�AȂ��M��D�"��\]��BsBN�xph}#�Z���%0J`Ѡy�ui9k���do��;���8����^�Jڊ|�3�;�����Ft�����!��i
��e_�[IO>o��,U��4�5 �A���n공ɷ�T.���ǎ�m��|Xƹ��@-��pܾ��<g��8h� $���rnZYjb
R6/j�hM\ag�{�Vd� ���յ:�
��?9��ʨQ=��A�V��2(��]�yW�u��邑 �8[a%2����^v`8s< �Rm�c*eYЮ�{VUģbwϼ�r��hLꇆ��S���l���T��h��i� !"qAtEN-�͐ɠm
�I6��%]w�o�>jg�~�K⁬���W�?~�!Ӭ�㫄��3+=��?@�	��ɏ��oD����aX!�?Lk� �Ajdٿ�H�69?�ƗG&��T�ߎ�mm1&iՂ�0)D�+]p^E&m�wh�6D3�J���ˮK���s}��I�Ӈ*]B����
̓T��FNkCW(��I��\͋)V�EKW��߂���A＇f�~dTl��:	<���i���mm{�L����f~����hĚ8�FN��^�(^ȝ�J5�5����!%J7��6j��yˈ ����c���Pз$���������1���!7���nU�=�j���xr���/��ߴ�H�?�L!�|�L��z�e}�忛�A�J�D�Kq�)c�FQ[�Y
f������O�`|T@���i���j���"����ؖ��^\Eަ��L�~� �<SΒk�!7z��Ǉ@l���ќ���>'�Rz�]��=�y³�a���q������i"#�u��*���*��>͚�ٟ)�� ��>��6�Q2ڪ`�:��l����Eo[�η��#������G�)�}�LN�W�I�t�t��@vî?@t�"!8ᓘc+Zh1	���e�7�.���4�� K��$��D}�C�յ�7gd�x�(�vi�,mTa/��KF\l��E_�ě��GR�Q�m#cb%�JA�ј���qsm1	ub9��%l���l]�������I�����{�d5z�eV������9nH/8�^�z?�~Q:~&]��l�Ã��5��RB8�K?�X������Ef�πY�kx?RB18�4��j7$V"��|*0��E�]
�� ���BI��@��g(��j��q}�����%��\�/��������ξ�P�ILH��g(�.� ]*��$��{����� ��I[�]���w}Y]B��b��w��nC,��;�Z����c�d�b �O��cU�|_�$�4C��/�@�x+6f}s�ĂW���YF��̀O�;�ر|���h4�_�?o8�������)�_Nm��:���ư�Z�`eS@q0�A�������!��doCm���#����wpt�K���n�D�/z��*As�' ���;�>S�-\%�W��� �5&�B$��Ҏ��:`W�Fܤ��9���Dޡ2�x)]1��MyaK�,Z�-K��g9>M٥ݟ�a @�ڈ�?���(�~5�a_v)}ߴo����-��}?jG�>#L��K��ej�܎�a��,���$�U�7���q�k�"�GQ� n^!�Ч��:�w4d]�o3Ѥ	E�E����ne%�6��۰��L��S5�d|��,q�z �%5g#�{�A�����X��S�*�����i�'v�un>>���N�w��C8藰��v'�!��\�|[]� �l�a����4ߣ3��K�[�$%�����iHJu�Ր�������mR�y��5~��p�Mia{��=Q�#d���I��g|*E(;X/�+M �S���4#T1L
8�օ�|�[�R��GBE�u�/@�X�HKG������5D�b����GA��޿"�����$�Rr�3}��˰ߜ�������,Ð *ԃ�k���Z=7 �r���i�ʌ�T&�W���-�͆�^@���+_3����'�It^t�ݥ2�������7���R�-7�r�	�K9����>h}�f=�Q �JB+ƤōK�0z�z"ߙ]���M���2-)�⅔�B�~U&��!�z{P#C�]9�UV�9ȣg�z%�_rVJ�5���w�դ��Y��g���~�&��_����N�99L<N��HB��2�����ER$(��]�p�\�(�'`�M��;6j��MZ_3�<�j�h��k�?�4md ���GK�=�wo\�4��sʸSj;DV"<�]����#����:�&�F��0�{�:W
�L�t��_���:�J�oL��*؃�́�Zoׂw���}X
9��'���b��h՚� Ͷ�kAw�w�u뻗R�f�S�nL�n�=�I������ȫOJZ��o�iz$�7l��y����|��e��G#��	���@:b��;��4��߫�'�ѥZ5!�V<��bMI���u��qAX轥�ڳ��m�k�-b4���Am*�<����m�-��Re�.$KZy�d���a3�n��������Q�-_I_Q�������VE�l$1Z(�]"ue��(� �kܓ�uE���z=�ωD�̖r
�����j�4l9L���\KGP�I�MB�U���o���9h*�c���ȩ�C{I߲1��4�6�V0��|�+�*F=��r��B'��'����aU��E��?�V������Sz ���ą~�1	xţ�o�4j�
���n��� K͹XlxVHYEB    fa00    1140R��F&��bܹ.�0W6^��U� [����Ƞu2k�KtG��o����ZR��墨�X֤�R\Y��F���◰�Y�6uAW��zP;�����a��&��mz����5E��q���a�!��Fe�����,69d��j�ǮQ6�m�`
�J��cK-eWL��$
#g��\�#�s�N�b�<���w�߀O$��gZ��'�M��W� V���ʀ���k��QHV�~�]�szn>c��?�q��c%�W=�;s^]e����ͰN4�h�?��l�y���~�������~P����t^�TQ�0ݑ��9�*�����z����9��N��8f������o*�nJL\M�/��%���(�e���ʟ6��N�PVjy�x���e�-.rĥ�*҆ ��)S��#�� ���)�©�#=m��C)��3~�^�����wHIw'p�S��4J����+��n��k
T�[��UP�
_����m}�	�ܾ�C<�ޘ�*�1�|�.�y_�ɘ~et��p�y��8T�����k�!6�����]@������8�n9�a֌�@�}����h �1���,))�eȪ�nY��rk%��`�%�;�g��25b"jn�\���[�|b���S�����gm�]�w��7������ǈ������1�����>&V���T~ʝŜ�ۚ�v�Q�vע���?\�M���=Ao�	�j�c��JE8���.AE�����=��l	�&���J�~�FG8D��ǝ"����[�|,��i�eǏ����^0��Ȫ'��/�3ڪ+�>G����xO�X����!��t}���ށbé�Gj{�MI?���Ga+]j�k�0IW�l�s^��I�*���
�r��m�Ȭ2K��`�?3�r;Z&���t	.��
��9
�Kg�� gPu!:4��Is<���5ff&A�{H�X����rȱSu�a�E�4��0�+"��{�~�%/OYn�M��ͻߍ�;۠W���E�K��3�2�M]�4��,�X����4#�$ϴQ��rw�ʦg��~o���o�-����Y�?��S=����Ӳaҡ�UKVw��Q����[O_l3E�⓴D����Vs�-@G������
��9B'��a��4�������V�!�՚��PVN�kxr�+����u��ӏ�?ˆ��r\wB �������i��ޡ ����9�Y�������@�6���;m�w��p_2�Xip̵k��Wn���c)5M��\�!s4M���eq�&)<�2`~�Ί�a5SR,��Q&3�z
^w���ĀU-mHD�������Y�M�,��5I~���h�9�$�b�:�P�rR�3@
���b���/
����}�@ޫz�e�+�Wy��͛�N����K̓�T��ܼ���e+Mx�u]L]��ɶ�Wb���{S�ۖ������E�|]�0y0�L⫱�꾏�b��u��Nw8�s�s��.§�7�ߍ<���r<T����;�o��29���#���u�7BS�����/ǉ&�� ���� ��<^��]�C��"y�~^��)9HS�a��%�뷍�*�w���w*��oX2H��AV��T-Sos(Lnи��R�tИ��p�� ,�����v9q�ޜ�,��J�/WL�J�Bb��ha�����be�ҪŪ��jӗ�ӆ��Y8�.�����ja�^ʏ1�:��!K��dWO��X:�_��Qd�D���kE���s���tF�ק6 ��Z��>�AA�Iҽ�ט�t0O��p})"Z�JD�/��WZh�[,o�X~WpL0Ks� �d�ƕ���,����aT����;�D�Te�Ly">j�-�k���֖ky��s4�ycF���.����9깜Q
�Yo�[���a_����O��>Z9���[K�y�@����!3��?ɢD�y��������@��}$�`S�,�ddC�w$IZ,ǊZPj@�Ə�D�1��7�l�|rB�������I4�v�?�lCq~���Y���k��"�Qׁz����3{"1�������d�5�p���lJ��m���I��=�V��JMX�u~C�a��t`q��S�d�O7�7.���:�:�F��=�[�G�ړ�d��aJ!�h�[���$����W��v:l
E����`$z��%��>�
�O;�GM�2�Sx�j �z�÷�!�$�H��ekߖ3B� ��cH�=��d�G�lJ=�Ū��L�({�wu�C�``d�7���2���ޕ�b�<�bD��<y�@��F�">�6�� 2��8,���4$�5cUR�b*b
�vqI�7Ш�G�1�n�9�f�B�.�&�0�wO��.i���ZJ�w�6�$س�Ɵ�1#�N�j��Ң���p����j)vh~�L`�u ����d���+��"Y1n��qC�zE<�H2X��N��VA��ԻG;wH��� 
63Z����%�w|�E�����Nh�|��eS_<"a	�˕l܄�@Iz�f�^"�F���A����BEg��։'_� ~g� #�P\�ko2���@@�4^�*Omݳ�Z����RE��Km�C()��q8LD�}�����ɟ"DKꗏ�B�"�]7�E�}|v)V~G5���.�"������ϥ�0낃����-QŸQUt"5��ػ�[O�:ܝ�p2u�����~,�K�v&2��,�$m�M�5H��ЬF�h��``ۣ��ϗ��R�q�o	�b��x��{�﯎��y��h�rQ�)��o̓6��V����+�	I51�m�Jb7���2��ʜ�� `c�Jm�M�u�
Wj6c9H
�ʵ�b��E)Xy��E��B��Ԉ��ϋeQ
�{.�Wm��t@h̃C�ժ�h���}����z�S,���Ĩ���rh9h�&�@fpR%g��=!a��í��H>��{�?0��(�d�&s+�Т�q��a��`ʷ���
��6ZP���'�bt�+�9�A��~+,�X�^�'�n�����	�Z��NQh�0�$s��Z�"�v����\xOқ��D�u/�e�T\�l��b=Y�Q����/�-��Ox�l�A����4d����
�����4햂��}��>�����"�M�^<fa����xZ�F��� 7�(i*}H_��{�N��4;O/�ܭBR���c����ÇK�=nqw�j���i����7���˝%���t�R~M$(��Ȃa,�&'>���֩O8[�T��:g�g!�����[~���>�l�U[y�[�V�iOQ�}�^8I�e�e�c�R���մ#׏F|I8�fI0K�k'�h �R3��+ �Aa��,s|�w\F(M�!����N � �ʯ_��3
��^�VCw���M���ZZbD�ZP�M5��w����%$jP��9H=�-�#h��G���P����Ž.�}֟�K%[0�Fऱ��.*��o�ɽlc'B�i�C���L�:��S�&2�%��^�q�"D�10��Ȑ7�\���ʻ�� �&�m v�[�g"S]匏!��`���ŗu[&Y_��L	�祕]�!�?6A	|Ű �3������L�-�dg2c����7����;;[��G�ĞՄm�p��c~���������Ge�ld�3�a[�}`�h�Vڀ�MN�Nai�Of��)=��B�Z�(�����U_̧�f�<Z*�,�
�������Y�]�֏e��#:Vʑؿz���݅��,����)�~RN�yi�
`<�R0�Ѝ��e����W[���� !ԏ�U|W����[�Ʈ��%����=����S���W���?{-�v������9�á�l��$T:.�ES��914�y.�����r��^A[�>����ڰU�_=V�+7�����7��,n�8��@��>.��;��Of�F��ia0���>���pf��f
�Z/D�D���rS֭��/Db�S�&�:c��{�YR%�d�k-�F�d�<��Ax���s4�^�9zyX=|��EO�!6�sFW�^�j�9���C�_5�0R�$!��:�����Q�P���B��=�;D\��>�[����y�a.�X��`��T�?�l=��E]�k�i���fk�<w]����
z�R��r�S`�#
�_�$��-���$�����@HAl�2p�fk��y2 ��N������Qj9�G�'��3��}zH�2ӬF���Il�E���[��ۡ�4	��"!Ш�����wG����V-��y����H�g��ᖃ	4�>�����y�4-�}�+Z!񹢵�5I�N2j�����܎yI�^g��*T۶(z&����+
_�I���<Z:.��N���I:�;��XlxVHYEB    fa00    12e0]&�W©q�F4w1RQQc��/�i��(�L�Bq���4����ǴrD�H�D[��-��l��4'��)�N��ۣ�r���O��٩)"��+�U�Y���N�/!���Q�`Z��w���w>�ȭ���^���3�j��BY�5ĵ���8�(c$Җ)�ꧥ�*�%?�Q�B��-��Ȓo���O������#��g�����1QC�1~�K�y�DMJ�	UY2�:c���YaӬ�7�IJ\�z�b�
u!� �g�ψ��6b�hv�����Ǩ ���~U����iI�
�L��c�GM�[y(g�����Ũ)Np�'�Bb�H�8^��=i.�VI�#��
+����%�(yx��_cQ�[����0ϥ1Y-���5����grG�v��a�5\Ė� �>J�� �zh��Co��!9U]��xHB�Q�L��	���Sb*��J�"x(��Svn��$�$1�T����2Ayrn���!E7&��_c��_����/!0df���c�c�͙�2�f�ѣ�$��]�Q�=����(��Q�V�g��X/�x��f�P$J�n<�Y~p6i�Bt���5��B�1t)�s�N�G필���!h	,��BD�����J7���K��¬u1Ϧa�� mKc�.l&ԑ�:.��(ʹ7�p�WQp�9�6��y7��7~vI�m{��x���D��Ve��1y�Cgxް֓��u��s2xQ��GQ$� �k�e��i/�I���O^�\�V��J�Ŵ.T�ݱ����rh�R
Cl"�s��؆���<a����n��2ɥ�튦�M	�Ibt�(`�j#�y/��\�Y�O:E�"2���*�OfW�☏盋��:s��u�� �!��#�.���x�Ƽ'�;���لM�7عi��lM'+`��N�a4I���`��QP�N��$;�%\���-��'ȁ㮚4���"{tLs�{���ʓ�+9���m��,�?q˛S)̄�m#�}��]h��{V��"��d%0Tȗ�
�e�Ѵ���ܥ��J�k��0~e)
z?�R��r�OXg�#^L��Ec:-VN�s��Unދ.���Um�rC��6y�Ko������O���R^�ј�+JF��a!e�v���������h�T�Ms��A��`�ww��bC�=z�{��d���O/�Z\+��a�%FqAa��?�;�F��H�hZ��\�9}0�@8"9&j���_���`Z
��U��z�s�-{ue�X!l[l��~�0���վ��I���|ɊFwq�^ǌӻ���d��7� 'm�V
R�0���k�,A\�VޖtW���i�P Ӧ �2���:��\,�]�Ox9D��ɦܡ��h�4e__i��j  #�;�
Mݕz���P��/*�"h���#OOZÊ�U��ɺ�f�$H���O&�c�^�( ������`I[-�;�bl��&���eZ���ɩ��C�ܑ��QʢXW�Gϰ�%5�{4����5�*���*�U��q��G�����.�9����S�6;���Ŋ+�P���qZh4�; �%��9Y@-ey[�נ�I��A�:Y�@h>�C�zy6�t6������������R���P擭T��e�e����FP���z|����%@t!C���%�gr��⤤�4z'��;v��?��^Xh�,m�)��)uf�C�E��g���@���)��3,�l��@6�`Q��D�i3���;k����(�fi��+��<��,�A>��FЛ����$��-m`��!�7�r$m�B��b�����k��tv�����ڹF�;��[�r����]�+z�S�3�O���?��!Z<F��ėr�� DL�|l�s�/��;�8P�xU��<�)�h�1i���܏� ��w����[Ѱ?>,~�N���s;墘���P�
�a>�'!.�Zu�x���_� s�g�Y��^��NOi�2.���z d����K��ݐ�,;Cp��#	]Q6eJ���ž:�!��b���X�ݕơ;\��,M��CAg�u�Ǧ���pK���9-Z��Y-��oo`��C���D�Ey�hY�����G+tE�?]����!���R�S���w¾�o��zu����AY%ܐ��o�B_-״c��7I��3q���_B���j�,*�4�*�1�����0]��U�ٺ��N&0��k�I�e�����o)!�2��,��ڢ9kr~�f���ǂ�&�Qc�t�ׁ=����!Q�_�Ψh��͜?w`#�����g�9X�9L�XRh%K��9���^\�V��G��x� ��IY*[���;)��t�Y�k�%��ŗu����d,�{�W��x�ȁ
S�
�i�S\o���}���]b�Y�#��0<�4́^�6�:���|e�Mö��[M�w�&�!��Y_!$�Aw.���+�g{�9�Xc��S�v~{BU��N/��O9ݿn>��5:ٓ�>�'�:z�@��jt�4T�Nj��S��'�w!��\ƴEcI�4 [C=�1f�$����Wx� q:q�*�����]�т�(��i�m����cj}���m�V���i�K�r�����s8���%�U����F[��9D��s�O���K��:v��.W]�4eɇLs��܆��P���3Dx-��g����&A)R�����
i��-,V���BM��˹|��t��t�	ޞ���	�w�ߣ�V/]#qXl^0,?�=�=o"�s�i�c����<Arҿפ�b�+j���3��N%�9�ba��T���A��U��j@S���N�;?h��� ��fŲ���5�E�Q�Yz���h�/@�%c~��U�_=�Lv��l�D,
�m���p-�Ds<R���Y��Ǆ�z�dg���Gd�{k�EjCAt��8m�G=��p+� �h\ٗ������`��Z/*I oU�Xg̊ǟ��Q�:�k�@�今�N�3Sp"_�����*��W:8�)w˄^4�T�4[3�ǁ86^b��2�x�H甜����c��lx.?-�������-H���,E�af��$��	Ȝ�T!���������̽j��O����i��|B��o���N����P'��_�~�#Tvb�'���{�n,������1j����2��ǌ��
�@e1��{�ת��]^{��H�����1�+�]�(EJ�(8�"[����q8nX��3F
�?l�Ch���5~�z 	�N��?;Z)�����<$zY%�1&~ox�f
<>�_�L�X�Y#Fw9���+����d^팗���,��`ZkK�@�U�̎s}d_%��k0ך=!epnmH�{@��Y���}�-yYp�$�8�V}!a�Qr�I,\��E��|��q�C���o5tkr�ݑ�X����N�u�֥I������ލ���T�K�~��]�5#B�An�����-8�6���yz扵U$��ljO�a=��V�ZK}|��?���s>��#��(֎���b��WENY��̯�"�`�ԢBrن>]�惣{����*o^�Lo�\n(�f�5�8}+�%0�9u�~%bvً�<����ʍ�J4P���������i�h�dF $�+Ԫ/I�z��~�G֭�������Pw�t��*�:Y�<;d��Q��O������qkݸ ��.�26�>�@��YU�,�[��V 텗�ƥ��cOH�����p�DeDZ��塅r�H�5��p�V�r�'�ف7+d���
D_�`r�(Bz��1d�3���s���
?UG��
H���p��B@F�Y�3�1��#e��Ηhs1��;��<�{��$�����|�r �S�:V��r��T�h�9�q|1��u�7�2qN�6:��?J�o�ж��/Bh�)��e�g2?�0!*֨�xC�J�~ 3�������N$��G_}(V�ha�v�E�H*�O%�9i�4���D1�,��H��5��U�^��YdsZ��0%URbf���+1+i�#�G��`���vr C��5�̟6r�7�{[gJ�]m�a˨���JoRi�_�U����4y07N UԢ8}�Eʙ���A�ayR+���_G�x���i֚���?��T �&��a�s�}p���,�=:(/uͶ���
 �?�O%9��T|���Es�	�L�6T:�&��M-ҿ��M�s�^�b3���\sD�a�X�\=�}	�T�[۫�8Q�ط��Kq��|{�c��)`���8@&B����J������Y����۔��J�_����m����-x�	��M_���c�V�w0���,B��׍���!gu�zb��Ĭ��(�c�$Q�mbxR����|�n�!cW�P���?#�'c�Tw���EŽFA҆�&���P�V|��}�N�.���Y�8�V'�O�^����,��r��U���C=����+�}Ȧ�X�5��=jG�>�Y�����li45:�g��Y�^�0M�>#w떹�p�s���+U�"�KĞ�ET
Ŀ|ra���Y D�/y��1X\���2��������h,���hE�.�Z6��8�6��Q�{��&~��?�O�=Q��{ouW�8��m�.�d�sTh�/S�G���Q"����������K׎���J�,C�{��4O��d}[���'�	q�Q��"Wa�.n�`)��'�ř8=��֝BP�r�\��`�a�Uۻ��!�)��WP'��[�i��ͩ��8����'�q�����H0�?�nC��#���\�g�	30f���b$�Q�6��W�?���Lw���gHl�Ư�x�XlxVHYEB    fa00     f50����Y�E�oqh�����3�}��Y�40���zW�Є��L�%���Io������5�6����]S��	l�ߒ�Dmm c6��P-�Dh6/1����U)Ѝ���/�K����L7`L+e%����:�k��l�9�q�5Et.�m�~��Y9�Ӣ��\��Gך%,~~�-m`�w�2t:�xcz�j�.{魹7�~�x)m�uF��J�z������t��e,� /HQ=C�4|�� ^���G����WF�v��
[�W"�V���tT&�W �5 ����>䦖�g&��{2jJ-�7�!)����˗B�(�!T�^�n����R��}�T�sm��ۤ:�gMG��i֩��ו�$s��� G;���ړ�pϕ���$0o����8ѩ�ܕ��"��h1.0�3:�ܪ��9*})��#���J���ʢ���y�w�,A`�"��dmM�� �x۫T������������Ωr*��:��[��|8,X�N4�&� �+�Y�=K�.��OY/�p��TȡWZ�O�x?:_Sg��E�������T�������^Mo߿Y�8R�����r�DjL��X9��Vo��h�!6AC��
�zԾ��GL�����8�{�4/�G��Mr��0uue?�-�d6�w!uj���9�/Tj�'lR�>\�	�����-u*�����0����3�Z���K,S#T��DV2髬�`N�V��&4��������za��Z'$�]�\��.��,,�r��Q�0�)���xX����mqÄ�>�[�^�g�B���t6v7L�dv��d��k��X��<?qSC�w�h�RM�y��Eٖ��R��<+e͗����?}�,�1��T'����bQ�w U��Vp:�.�����X�:�U���1^~hQ�lO���)r���Ͳ��6�r��>�
-�����0YK�!��>���Y�UZ���m������63�3W�X��?$n�]�5M+��	�x��.�2��� �*cm�[��6��~��)����D�xx�C�9翿�@1Jo�&�^�s�uM�t�{ADqF�|E	&:��uχ#U�a�q��#���V;Q�"��@�CAb͢�g�����"���r�??~�m�������[�,��h�4pP���ra�D0���Y��Rpa8ڭ�a$}7�-'�9�I�O�OVD ���tN��m��Y�]k��Ɯ�Prw�둢 ��n�C*�+�V���_2� �-S)��X�Z�%�#��q��M2����=D���-�q&Y�Q�C6�4;��2��wdz��xډl�A�Y�����ꚥY�����D���Aaq��AUD���lE/��G�(���ey���YW��H-�z����0)m6���#�j��wl���_L�s|�i�4PN��<X\,����^OSg�8٧G�E�H��?��cH�}��A��'+����9���*~&b�n���	C!KIx�Ü�|�(�愹�_*�r���aP��bQ�+���"�^N.?j���d��)8a>�q���\�_j:v��Y�K
86Kh>!�����aG!�ƥ�jK�T�����D����g�|���j�K]á�{dO"	�t1�����&��y�,m���Z����Ƿs�g����"�����[I%�} [�c@J�[�|�jP��f$�at`�������+�x?�C�ֿ#E�|��yN!�:ẍ���U����[(4��C7R�>�WZ�+�Z#r�5�A",�!ꂽ�r����L��$�	�q�\�0˧�N�j���*����! ����2LN;+w�xF쨞�H{fwÔԟ�|��G�T�cO�e��kjo� Pޫ�m�.H~�f ��M���nݣ����>���8�T6�w�w��O����} �A�d��pI����|����MJ�N�4(xE���yM$��>A���?�bN�W^��T��P;��jN�����5zv�W��]�����m��.S����u^V]�x]�7��oZ��m�5L'��Q�"\T���`Ĳ%��o ��L����sgP|/HM�ё)D�����9���8�I52H����HZmĄ=.�j:�?�z��qoDje�R��٤��96+J��������w���+'x�Uā_4z�_u1���[�i�-�b&�6�s3fY���?��*�S�3EA2�Q�u�L�pW$�� �nE0��������O}h���榉�������E��F̹�(c�X�����%�	��ݐj�[����}����^����"W��R�62a`^ 4f
��'�g�F4��]����#Ō�:��yTa�g���������QCtwYl�7 �[�4���&hC�y��S�~�y�ٚh�����=~��Ec��0�ڍ�$�.CEv�
�����{��g]>y�1u>X����\(���R �T���N���x�T�1��Hq�����$腎���t�"T��t+��%�����=�YKCăG�#�,}t,_��D�KWsKd�z��u����K ���~Ic$L�~�wu�*a:���&��YPg�a*K��A���\��ZX4�R��#ud����@.��)�R�L(j��{@.z`��o��,ܭ�bijw8
e1
�y�����^�
#�nz��'j�/|4��0� FII/�N���7����OpPy�fLzA=��Zh_�PlB8��'��&'ܦ<�?��K��-�:�6f��#�k�ϟ�]X���37\r����<Au9c��P�d�lf��%юK�k�Ҽ][�z�"�hZ����C�ׂ���V���",Ĵt�9��o��G�C�]9�V=r��؄��B#'l��͈��@�Y-���w�0�h�	Iw��$Cي�e'�����v0�tY.7���}�tc��_�q��e��	a��#�K���F����>��P���JK5��U�[�F�%˧K�-|����{,H�;��Ja������8�ۓ3��,E���|N�<���?��8d�Y?�����g�u��p�7�M��H���~��ы���F��UD�_2��3�4
.?Ӗe�P~��\�E�"��[�"�9��OA����	�T�-���A��K�]�gj	u�zfA��	�0"���%[{�D&��m$,�����Ta���/���1b�QI��߇ �r��I�M5T�#��i�TI��%�xe�t��4令&���~�߶5�R܊��^n�g������|�`�~�M�=�u�Z�坦z:�Xd��f,����}%���W���L���{�ƇL,��UH?F�vk�>�����U6�H]}��$?V�����	ב�hnjJ�n�t }�krA�hۉo�q\��cJ�� 0�6GF5 Ƨ�f�"�D.�v�myL��Њ5W��٤�~Z�|�*w���nb�D?� ��u��3K<�Ѳ�oՋ�*՞F�ȫC�z���zY������]��s�O �1���.^(�݋	;W!���!�&~�,�&^z�?��b��7HgU3
�N�P���rAT�PE\C�_@KU���8��@��1��z$�jҕ��Բkk�I�s�����I	ʣE�j�TRF��I�%+fZ���&�S`rR-l�A����ߣp*F�J��(���� ���v8��)e>����;Ag��~�c�䑙��Ht�6J<
B:ϝn Ày����s1k�!/ң��������8��-ԏ�һ��|��^<����������d��Mހ�8nr��Aw�)��*>��<O��O�䅿�L�[x!�Hh4]����?A�AW�}�L�,���������3TU�����̻	@������j�Gj�l	9�Ev<_�!���;mC�גP����:�_�f$�ΛXlxVHYEB    7273     5608F:�7*n�I�H���u�-"�B52��j����{M���[�3[[�0��~��V�z1��(���;����O^߬���g��t�*}��)?�����WX������urF�45	�<�1f�3���6m�4��v����)��Q���v���1��2��Z�����D4�2����Yǚ�N���x�'g�tՅ�Kﶱ��#��$]�YE�)P@�!��c�:��g������^^�����E*�z!df���W3�@Qu�dt�UPُ�>�������vXZ�Q#��5�������#�H�3���	��U���,ō<�j9�`����S�W�jG�J��$:z$"�d�ɷO-M�6L��a�B�c��n1��F|������� o�{}�4석��]�CH@�`@���J�AۇL��(׾�`������f���ûU�����g��&�,�������"��;����m�pq!�'z`�ȓI���b�L��/���OEP�Ϟ���)j�;��>��YJ8U�X �֜�#��� 1������h�p�Ė�8��Ba��<(6�r�z"!z'�fa��M��~�g��}�⯦E�^To����#�m5~w��v��#�|-�k��qou��jU�XE4�A��}�P]���#���?H���o��?^=�Fp���3`���~3>���gpkA�3��Ҥƹ��w3X�K1����0<�%e �V�7���E��9|.�.ڴB��,0����1��y��V3�.�j�&�QV��>�풌m֟�
� _�O�y���\c,J﵃�^��$�Ky�<�������Fx�v�����a>�xPt����~#V8���O^�_�<�/�x�%�2�Yԟll���p��h��`�B˖t�Dn��6�^\�����l��I��YH�O~j��Wԥ(��CN���}����QvK�ӎ���}�sэ)�J1m_V���ǐ��5�QN�3�պ���ے+QQXP!g�O�? �)����~�"�0o�Z�=̧��%7���M����nI��
!�9�l)wn'I�����J���}�W�v��H�^�q����݀9���'I~�K��cBH���K��� �S��d~oIsJ��?o�,��
0M�e��+o��2"Ī�ܱ*����c����� �{�蠔�#
1{��5���'r2��`si�3^�GU�(�V�6�X�=q�¾�{�C4J�A��w��݂�f�;pM�I� <��7�������+�ZG'����rqCs���fʝ�2{r���$3JS��	�{�~@7�HP��N�V'�ɔ�6��+wWaҜv�b������:[�l��c�jN"��	���k|�i��'F�<r�ܲ��