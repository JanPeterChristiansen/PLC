XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��M���A_��?l;w،[oxt
�T�[�R�Wb�J�����|+k<����f9P*�T����` ±4_7���#�"�3$:�����B���/�8�\}��`8T��>a�	��],��ན2���r�U�1)�2'b%*C�6���#���;�k�����0�Z|WX��֧��ԅ��C2.rkq ~�X� ؓޕza(��y��ͽ�,�	��#r�D������f��)��?"S��4�/���"*� �8:��Dux��Y,�_���?�l�$��6l��}dA*H��MYL�[O�a7� e�ru'�ENm��m@����8iu�]�1���ITz�������9�~X�@��/�m��}c��곂o��F-�;��D���r�3<���;��u��8�Q7 �������K
�ۆ�')�xaw�*����n\��� �7��Ǐ�5��Z�Tt0�
�@b��ܚ���7m��,��TOz�E�^}�b���V��끮6���b�>WFbSb�Mm�$џ3UѲQ�,%�5����������Ej��<�����Y@���!%Z�}Y$[��]bEA׊�OU�±@Ac*#��rNk�VZԑ�{0��[t���ztfW��!��x]8�Ʌ��2���i!'�egVp�eYʴn����7L��r�G��h��-տB.o�P�q~	A�z;��9c����hUd}~��0/����N.*���YH��?>�$��
�&T/��k�6m�T���-��_Xff����XlxVHYEB    33bd     c90d  _���n�+^د-�3ҿ�|�y��P..� c�S#�(���T�pS���h��Bh���KWo�ƹQ�}��r��G�=r	h�:R���DT�&$��m�tz��ￌ
��)gOi��d������]Z͠�a�l����=���Q`@��癅�KB�����;7¤P�X�����/�DO­�� >l5ܜ�X���~���) �󦲯���^�Dӻq�w����(��"
���`��j���-(L9з�[��ݕ��H�	��|�����:�զAW�SN3����.ުc�{�B4U�z��?�@!=�>̿X
r�2?��Q��1|�>�g�Zg�Ն��d�}��k�m[�MCE��l�md6����v앻+�9 #�+�i�n߭Q)�����ʽ0W��=�?")g�@=���}^�/^�>�G��o6��4��*� �`u<�m�`��ʲ\$��f�:����r�� �1B��Ǭ��A�&���x��C_�o��~ ����@�g�K'VÒ�4<�;�v�8�#��6pu��1��_�8�����~h�lm��;�7p�t}0jw�h�������C�ƛ��/�rdO�]k~�p/�,R�����y��c�[�=�7�Sa���6����Kkk ȕx�[�I�2�c����.���t����9��	��y��d�n!�cR��qN"ql��H̱�t�8T�'T�:;���N���&��ȗ��sT����$!~;��C�(A���E]���|!gH=��&��{S[_
3F�Ӝ�K����Ӑ]���۫��c5�ݜ�V�z�$��;s{'cP8Z�@������
��7o�֑�ƒ�j��E'T��D������bQ(���u`}�W�j9VJ��Tվg����8���8��b�u�W!�̦�au�S��s�ez�d���Mr��O����IJ�凧p�O+ƈ��[
3�\��81��hѥ�&6��.Bx+���הޞKȋk�[�:
�Pz|Lo�}�|����MkS��e3]�����Q-����@<�4b�2�.{�=d�Bj�5�9��芌�lTDO�Z)��O9���4�SEԅ�����ㆢ-��2z�#SO�t�x������{Bٍ�8�����6��D��g��q����� 4fޔ6H�gpK�o(�O�Je�t�횸p�7:~×�I
`MP�ө��)2o�8D|�����q�q&���sS�)LY�u�s�]��@���y?�Gu ���R;������~5LJA$)�� )5�fe�v�+�����ߪ<ʞl���~F�0p��0K����<@o˖z?ϞK�wE<6r.`9�����k���к�=Ěd"�{�����r$i�\���!�$��t�9D��>����'��vw��$��4Y�CY�it����Ê���]A�%e�wy?`6�d��C"��u���E�=m�ْ�tK|l4m�`����`�S{�՛RA4r���c��7��$@A	�΄@F�ʡ[���(�6�8F���@r�Q'>�
m��v�6������|UJ.�īK
�6
U9�hR�*_�����p���pa���z�jK4" ���
��Sb:W
��p��Ԙ�R�x�`��p?�g��&�\��z�~��nQ�3>+�J����oY�`�mg±0�ʵ���ؐ�P�p�r$~��_""}'����_��}Nm��oT���w��k��к:��Ŷ~�7�6���5nP�N�-��;�]�u5VIb�hf����>ڨ�С�$Y.;Xp��9���a��h��(v<̟s	�XN�]�`}0����&�#�N��z���>w���| 5�U�	���w6H2mӵ��5U^��g��~GI�˞���k�K��Ck"���~ �k�$���˴����z?�r���xL�����/I�$)�w�jR�|j�]�]v��݉-i~)���ʡ�P��ne��#�OS�ˆ�32fYQ&LP�y�{Dgj�� ��J~<���ڲ�?��P$ѱ#;��� ��}��
8�^~����W͢O>�H!�Q�� �UŴTϊ���
Q��U�tg�M����>&��1�}�+�܋v��or�D?���x��JHL��8
�U�K(�l]]��VP��4_�h�*�~MKW�M�-ܕD, �/��NU,��P ?��`k{�Ns9)�CM��ٚM�أ#�l[	��-?�<��p`E���3��ᗄ=L����g|����\4�9�:��LI��.�	�V�l �Nw ���y��s�Ǻ,��էm]"�7�F�78J�J���7t��F7�d����o��i�����NͰ�G�!�qJ�n��Rmh\�o�3O�"r#8UU�Wi�DV�J¥
���#ٌ���c�΢�O	�^��ë�:|H���t%���1����'UvL�ҭv62�V�J�r�r��ȡN��v������Q5F����u3��X�޾�.q�,���d>Ҁ�s4>v&y*�� P���C�IzF�W���#ݥ���[�������X��b��<:�l����ү�+���g�lO?~�9|9��[�u��S���?�XB� ��1LL���~��]���K���v��1�2 H�!lG�C����͓_@̔9/G��⹹�Ʋ P�Ui�
n�rFѡ�I@�eύ����{4�ë�Ґ���D2�*bm^^$*/���xF� ��] �Y�O��D �T���B�Q��J{�\���� U�z�bK;v�a�#�b�c0l}����P�j���oY��9�D8��(q�i���۪O�3���~�2����p�o6����6hN=�k�����l����ھ�k���L��zط�wV�@\�&��5
�i��o�`Z�&q$�#Xn8�Q&�>GN�a��Y�s�8�7b�'2�N~&�IW|��JaXT���=rv�ȁ֮/Pγ[�P��d���x���#ߠ��Y|-��L�T�L�� ݒ�;��z��X��0���(һ�p�+��(�>����*��wO�]�UT܉.f}��.R@�%*v�����Ә��.�ԛaL�o"�t�; ��C5ju�hu�H\7kSZH6�G���;��=�%��Îs��d���Cj�e���ϐx���N:%!�h����!ٶ�������v�3]��Ç���g�|%�@���