XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��:�R�3��ؠ�^�����V�z�R9�4*��5�����J郥��2dv�o�����c2��&�s��������}��<�f�C�싦��)ğ�y� ����j�l�c�u������e���WTU\ޭH:GW(塇��X�'k��f�$�yg�� _��޹��?�N_�	XU�U��	���L`B��;7e��QL57!�=��f�y���U@�«]
�֨��E���n'.�{�D�ϱ�9
���(��D�ȇv�< ��mp_����d��h�R�j���0�#o]
�K�$�:��Kڂ3���L��윚�=S�l��BdD��q�B�Ǹ#�b&��>�}��t��	0�"]e��El�i:`�8MzY�Nz#E>��^���~���&�]��)��u�������"��IY���i�c0OL�V��P`�#7(2Ti��o��v��%�枨����mU\��l��������_#������
��I2p<Kq������J'�O�F���1��G+/}���Y�D�3f��F���E�-�l4�Γ�aMyfS��`����:�5�Kk�S���E��>&U��4��3��U��u�'��x��`܌>�vp!���+��{)�@����~G[���0âoyH)��8������_$���Д7��@��$I,55h�H�a1<�P@����H���㿘W2�z��] W�
A���l�h�B�����%u�9� �א�P�um5�OZl��c�q��L�9����XlxVHYEB    aa52    13d0)P��L֠6ד!�/w�v�l2U�]\V.�"u!u z��V��C��e_F��*�Z��\�-��-運���'�ة���k�}V���Ui�^ؿQP����� �)�-� _�*^�p|�
��괚�] �Y�ds��&��0�n3=�@p�v������H6�o� j�(��ꆸ�	?�x�h�:@6.���u��F2�{� ���Pn1֙���U�&ט�WR0�9&�P׏�DF~*�+�W�"���n���s��R�"n�s����/���,��W�Zz@�I����]��W��Տ�}vK'���N���1UЌ�Y�zU���!�j����F����Y	�F�Q ���i��`�2����q�ȅ��m��{!�sa�v��)mR���\�8���F�PX�;ql�̺�V5���vR�W2D�J�lQ��#��p�]�����]ntL)����#-�W�����/>��H����q�p�D9��������@�'0�c�(�H�������M ��Z�0��7t	�_� j_���1�@����s��Я�@	��G-Uw"|kz}�����ӓ�g.q�ݏ��b�޺������ꪍ�@�w�W��`7�|��_y(���\�C
��
T@��o�O��ކ�1֮H���t�s�JPD|6���X��'�W�(p� �����1몄h�cפ�,t.��~=�w� ����>!�)KS��a�Y%��ɘ�~g����<?����-h�{.��y����Χ� �̰X]�zHv48�����2��=���{@~̖̭���K�{D,c�/��)u,�pǡέ�c	��!��Yyo�����]�W�lS2��ޫ>
Ml�JG�1��3��/����Yz;]��+re�v@��!����xl�B��F�� ��� }���PɁ��ً �� lh�5� lE�
]��.l�@���?���ۯ[u���@��DU|��:�����x�)�+��!�t�ԤF:��C�CҚ���C>zyN��$�V��������F�T:[z�`lϣ!�@�NXm#�o��f�6�R\BZ�����k
!��N^�TgRad,����/	�mє&>ܢCvCi�}sM��7�ڹ°}4�<;��i�P�Z���n��nO�Ss�0@M^��Q��Ϗ���~�bV�����ԍ(��9�����A�"Z��t}���R��5�i���80q����αJ�@Y��� ��Axb�D�0��g���l]�j-�C#���e�Y�8�<�Ijp���q+�f�jX)�������*�FO�f�ݸ�W��Cn�N���d?�'����g�h� �9��5Ε|ig�$�:�m����pU/;����9)��#_��L6�d��z靤�ѸX�\��btϫ�W�y�gUIߥ�P�Hm�� �5i��Yg�$�z���'�5��D�|� ,�|���g����F�Ԟ[�KU�V=Og�>��=�M�T.�Oy��Ӈ������GV�S4�����O��WgS�~��_������sk2����N�p�(��DR�K��[��͘;�,����I���Au�EV/�E�0Jld$��+f��Ta�H���������w�W�oґh!�+ַz�$j���|��*�3y)x%�]�e@r���+�핛Ԁ�sՇѻ ��됤}�E`��"4]�$����l��F��A�q�Fi�D�0�]�̡hQ|���k�6�$�4�!��Λ��:9T�~��,y�Z?g;)��Ԣ��GZ��ߒ�u,��ҹń:�ak�^�bcA�цX�Z={$5�l�C��j���T:��~���eE�N~V�;mY�l;�f&�k�б�K�7�����L��i���)M�"����O���1w��=��{�,-n�T�ޫܙ!@u�mŪ��mrPif䨯yt���%@�\�y�)P�a��m��j��k��@��;44P�u|��D!��l�)D���G�}�yצ�]j���m8�z��u��V����?�-�4�s����3���bQlR�Cu�d��E�nž�+^d��<���sC���&Lޓ���j<�|G�q+c��Kv)$G��v�����sO)�(�597��C�''���bWw�T�^�����5�j;�F7��H �Z�/]���뛅�%]���}S�+V��k��͑9���X+�@4�OǑ��ݶI(oe`�_�_'x�\ ��>��3)�T��W1	���D@8���&�ܽJ���3oK�bDi�ѳ�2�����z%��C�h�3�2li�h��L����������#��?��ă�@������bR�Z���ے4t��F)މ�j���>��`��<�Uc��^`HɏZ��q�"��Ý�{���(C+GK�@&x� ����Q��:�J��>�g)2����R��q�(W[��P: �~��%����)��z/��]���zy�R�{��1�Ouo�v-4&b�/�)�2Ie���፡�V�0���g�Ziҵ!e1�kA��2l�M�R�l�ih����~;���KB�$�@W��ՖxZ����������m.%�a��H�� �R̿��`�Y�$��͖�2lim�&&v�r�I@�Nq`��	t��
�S�}��Qϟ�5C��mH�Y��g!d�����)O$�0�\mb�
0�zi�\�yUw�[SZa�|0	���3�U�Q3��t���������^%�*�n���:�l�{��Q�=�A�r�L)��6^�
�0���r��$M��9jKX�1s��sTF�ж� ��&�ԧ^�LG�Vye�KzM9"������#�������@tC4���:����2kol΢�5%����R?`�]q��r�%cQ]{2������줥����v�Иf��$b�3̋�s�`�D������Ek(q$�Ag���ф�y7�!�&�2_1��J(�>4u�fC�b���RZ4�b�,�
SQ����|�[P��)=�0{��au�49Cت�����&P�K�F������(�Ka��d�]2��
��fL����ދ��[��xrW!�i���J��	!��Kp,�+����{H�V��S�����q#�@=�۱�Ԝ�W1J���M\�1�{�kĪ��{s02��������dI$��lzP��bE��v'˸-�� ���d��.�}�_r��J��s:�He�Ϡ�d��C�^n�:q�������vύ�aUr�А�^rk���R"8�e�dLp����.*�A@P���?5���V�@���rE����&n����.��,��=~-L�޵z�27�����'��q|�]��Ƀ'uw����IW�s��>�ִH���/D\Pmަ���#�)�֗8�C�ػe���
t��ȰDxz�ˇ۟_�)l��PϬՄ��#�8�WbQ�v�I4��/��_��C0o�~,&�(jf���[�1cx"gC��o��h�3���X���I"�v=�dϪ����E�SP}2e����+ګ:M�<p�&ѣ�Y�,���f��>>מ=ce+{A@՘��@d,������y�A�Β@��4YFBnHV�`MWt��pc�k������`1�*�����#�8����miL�$���e�7��Ӵ�d�gHZ$�ǂ(H�וE����*51n��J�"Dk�]c�l�`$zqi���+j�K��XN���lR#�u���uHꛘ�O߭���{Hb]K�;V���0����T��;}�7S�&�mp<�[tvm���¶\̃����J͐�����lh:�c�ۿ??�a&x������?L���=7�Wj����5���b��|6 ������l����W"�*�!H�Prɜ�9R�^2p/[g�~Lj�d�	˜.��)�`���Tnv�6L�*呱F��T��O�k\���իGm���o؎/xz��-�=Cڠ�K��e�](P靑M!	EU��e͗4fe���p|����k��tY�?�=uʣ�L���#�U��:���ZG���M)�o��|:Se授V��c��}�4��Ď�{�8���٬Jp~�
�}.��sC�Lm�����Q*��+��x޴�a��h#�Q�;�~�����ؼAH)�Ի�\�̋#]�����u�;���Zfn2=<�n��,K��w6$[c��8��C?~�t%�Um�s��Gޤde�b?���ǬL닱S���ux� uO��XQ�@0�8�m��E��}T�ԪV�ǲ
����s�K��EA�\^r�;���P�W����m�B����1���.K�G��R��n���;�N�����"�,k5Mv�_�-m��G;0b���Q8�|X�pDa�o�����=v�n�vvω���F�,+ %K,Y��X�W[5{�@}A�Ыe˚ri�q5�P�:!q=��{f�~��K��@iLҖ�^���y�x}pĴ���c�k����Qj�3rw ����� 0(���I��=���5]�ea����|��@�b��쏌�B>�ˌ�`,��Oy1�?~� �>�3C�w�8
�1�X��]f+��rz^����uO�R#hU��E�y*�Q�\؀�=����F����?;��������*́0��[�����t�o#z���Q���|e�O��WgA)�,\��T(rn��C�(]�3�]�F��Hi5�d���25liD�!���/f�MS�Kr����|��U� ���;��]��,L�7$��}D�'�zO>�z02��v>O�lܙNc�(i���i�x�n�R��G;�N9�cSe���*!�"]M�hݪ�I�b�G5(�&]�����+Eo���[�|b�I�|$0��2)�e�؝f��a�P��[nO�{�#�+�]�6���\�������u�z�d��ې}��y91��~,"n.Y�C��:���~y�JS����Y�Ƀ\S+.u����(��