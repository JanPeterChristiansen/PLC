XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��;�-!n�N�RɽZ�x)�Y�(:�=_MJAh��l���C1���׃�����x�[�:SwCO�8�}�3OCt��8B�t�XUO�K�i����U9��G�A���њM�6h]Cqb]r���;<Ne��,4���9�_O#�]Z�:��Tr���O�c-�-�u�*4n��$��F T<��T6q΍6�_ս�f� 13�;��X�}(�����E�������д����3�dƵ�@"�ʠD��B�h�6���j���"��˽��F�|t;�.�Y�<����︟y��O"��H��C�Xl_�p<��r1�p�j-��'��#�Fx�7�g9�P����N����FG[��h���=E�\�c�����V�**�' l��@Y���,A�����	�[Q�k��R��H�r�'p��0���w���,��+�ҿ�>݋d�X���b/�[v�e��� ����S?
m;q[�=����2P�����"V�N�۲ ��H�L��� L<h�9	v�n��)&v\��{^��� oQS8�>�����ܯ=[�t��%�{�c�5gm�Rq�W�D�̃�����T�Y�&D��Z������0�������Ϯ��ꖮ,�z���.����]Ji�{����X�A�p!�!b���Gu��6�vk&˗�����R�˟��+I���w��m[���w�w�"Ŋ���n��l9��J����gp���Ý����� ~����͌�XlxVHYEB    b631    1a00*ܑ 9vY^Փt�<'��Ԃ!oݹp9��bW���;Vٽ���u�����$��F�کW~A���7��=E�}9�I�k>
�0sj�z�_��[����*�daa'n���o�)�S���6+#W�r���0�M�"NI�����*��>��氹Ϲ�
�w2y
F\�?��(dts+>��SlQ:r@����<���J�������r}�F�:��f�0�t�n�#�@���m%ʪ�P�~�
0E.xXZ�|���D��)��� ���W5����X.���چ���t��k����䞎G:�J����p��c��k��\;%7�ĥ�Z����-��7X[��K�S�����e�J2/8cv�����H'Dh�-L� �o���x��Ԛ�sTG5��9(�W�؏�%bp��Ȉ�)6�6�dO ����/3�?�Q�j���)�߿��Nl����r�7�*_����\���d�x�����IW>��Mjȋ)>J���(Ǩ�����<T-�����?��̦� �r��eQ})�*�����KcRS@$��*Lg�?�@���FܕH�$��\)���1�!V	9�^}V�T�9L �� ��^=�@�HܨNNzݸ6�A P����8l��0��Hϻ>�O|�D�{���D��3���ˊ3�F�;mo/Ih狮���ub������>�s�7p	��/ͦ�a��kdk�>>k�N���1Z0-�,	 ]��q�=@�Ρ?�V3���78���ʺ"�кc��(�RH��B�W1�xx�	h�ty�5�����"�:xo��;$x�A壮<�M����,���f���~����<q��nN���d��z���� 1�)�z�WqHR�-�úNn
�x��f�p�a�B��d������R� �hETi3�J�������k���� �������x�#D���0���х��݉��Y������b�ʻō9���� ��d҂�';�{�˕y�9cW��8���E�0�R�}���D�i����;��9�۳T��u��]��Fn�?�����sO�Zl���_3�0t�y�=��h�H=�b�ŗ�U��������[�2$J�DЖ��|%��P��4���u9;��|;�)7�?�*h��!St�>�Ll5�dʗf ��3{���nw�2�qǕ���h�%�&�����K�S�v-��xXp��_��
��A��F>�%c�
�Y���� 0с3���ܯ�߱����H�� ���I�m顁L�FN�����'�w/����8F��m�mȸ�<�`�'��`?����E�S�P��Ӥ�Ĵ���Bb)����BE4T D4�̯�9z���T����w�n��QT�"yl�&�^Y̢�<{<c������x�7b���O4����T옸	�y��l)@��SV>Z9�O�%ͬ�ᏄW�y2/�`՟�,�FA��a�Ț(j����j� ����%�1�@ 윓�n������0�Ug�������5�+�F�c��w�(}(4TP�F�yJ}���X/ ��0�f��v��7�^1���u
҉��S�[�f��ӹ��C"gi�fR��D^dS"LQP��B������.z-���P��^�Zo����¿ߞ����2<i�C����8x�nN�6�0����	��.���OƐMHS��R�z��X?�+N�Qf�>�\�����!赥���p('�܆�]�f���zRb���A�d 9��.�ks{v;��G9`3Ο�n�$�[;�[�PV�kr��Qۊ�c�ri���db���g��m�6��S�T���H?"=�D����2����6��`��q���}�~�P�h����=�U)}ˇ��=�C�~��� R_b+g�̑��(e;z)�(f��X�6ι��T-`X�,�'T��\�ܱ��s����pf���ͽn�!�GL��x�@rOA�/����<�Ņq4sa4t�x��B��K3k2VE?j�Cr��_��� "g��OLF��spo�W���T����#��s��!��Fz+:������;�%����J�zLb;�Og�^O<�Q��2�6~�ڒ�
Ow��chTP��T�8����i�1�wT��aP�aI�����P��;겱� �K���s�����Y����g6�̰�Z6�c���$c-��� ��'�^R���qZ�ܚC�o�Ux�t�ui}3����X\����}�
p�K6u���e���#Od�ۣ�31`m���K��L����Z���c��@{s&�W��sD)w��:E	I����H�bc%u8�$�1KѠ��:I�UZ�&^�c�w�ר�4j}9S/Hf�b�N]�Y���_V��BAE��˶�cgBݭ*��SGr��I1u�B]|�j��e�8��*_9�u�A��������qsY|3����ٲ������ٛ��0Cv��9GpRx��g�SG
_BA�Ծ����F��l��'���(� ���B���!y�h�՞J���P�D��t=�#�%]R@i�N̽h���������/�v߄����y���yp�� ���,R�>�(�m�L2c����Uӛ��}"<���T�K��2�wJ"9��P#��`�����u$�[⦧���#���t�(йAĆE����'�rh� bL���~��X.	R�lN2�
����bj\�em/c���M_�T�/r�u���d�ǩQ���}y��8�s�E���;A<�P�T��X �_�s#]}@�e��8&)㮟p�}��O��� JY��g��44� ��2��g�#���D^��8(�ƌW)�S<��X�)��Vu��� ����B���"L.���K��+$'�e�- �'�i$�2��@ب���#���K�'�K_����=�q˳�1_>z}G�\�gWZ��� ŚH�w�'���|��ԒZ� '����׮���̮Zt�l٣<d�8���Z|�EZc�	��xG��x�ϖq\cBZG�Qߖl���tw��)Be�10X��ƴ3b(�*��dY.��^�(4�Hh�ɩ��)s���囹�O���_��PxN��4k>�H�R}$.�ǔ�݆�|r��v�s$u;�#��&C�r��UG�2ry��L_��j!���4���,L-���ނ��
3�=e��:���pp��W��xP�C�o��I~�����]�s�\ѸE�sm¿������+R�(mx����b�;B�O@�~F�ƞ7=wCK5�7�W��y(�G��z]֎X�[�D�X��%�腧D.|��G���RBW��(���fyp�<�,v�qn���,x�8#��} �^�o��k�xA!h���(-갉��b���_��u
9��VDц��ĳ����3�"0˼� w����2��� ҭ��{�;ʄV��;�bˌ{�6LF�L4�|x�ܹ�����ؐm�ڨk�@[Ne��О�{ƚ0�n!�����nY��R?��|;�#����.ʙ Bv�����T�
o�c?���X��r)��d;��[��Z7�஀�s�Ś�m�� 	z&�%/S]3i��i�x&�M��SE�=;S���d@L�|]��oo[����!M:��m[��箟�����crj]'�;����㢕�,��)<g��+�!����n�$Q�K���F(��)�;ΐ��� WJW��4=� xV�fE{(�u�V5��v mޭ��Czh�&q�6��U�D�	�o<�lDD�q��c��.�-���ן�|��s@�2Y@䈾�0�d|��4d��L���Ըse�o�ɗ#@���y]po1u�1\�4��^�'>�v䋼��<Ur��d8�k{�s�,�����X���U��
�cR��Z�Ys[܈{ ��s+�>��$k��sv��;v(/���`R�� �5�q]�8�o�
R��N�M3�t��h��M�oNC uk�v��ȶmk�u�����x�>z��7�t�G]qz�<�؀����'�v�����` w}�+�T�||�]�����[��}������~��QN�7���̛ɇLaj�RJ�Ɛl�@�5�oPm����S���_�7���{�^9�M���9��6�+�uNn��8�S�(3X��E���M��jK��F�2�'u��Ӽ	o"k��e�L8
�����D��_�����-g��:z�l+���7ݗBL�Srg��t�U� /k�o��k�D�IM���G���Su����|�-�~4��X�l�>%s%O0l��i�?��e#���lK"�L��x�ߚlj��l�
�@�L�1�O!��p�H%L�=�E��^�moT���SP�<��8S�Z�5�����d֏0�Q�_ �����k�/*���0�.�N��5[r~�:`;��KR�u����/�`U�2�E�2%n�~��,$�("A��)��m�ÐS�XC���&a�1Df��*|�D=0�d�%��V�^� Fo�R�>gT���r�iD�S�G=��_��ݟ��J�Gk��
gp[�$��Q�Ж�~g�.A��åtW*�K��w���ߢ������w�+��~��q*����ZϚ�q~u��d��FG}���W�a�D����Ĥ��!*��C�I>'�C�$p�ŵ������jh��=t��?�*0�^^���ޠAQ�_�_e�&����Y�E#<��������=���; �N\K�8��fgA�y���;�����&�S�*�'����0��B�_͉�>E�ޱ�<�m��Q��3�Q5�*�s,�
	�J�P~���ᭀ;��{�[���[=G�|ܓ<�+>R�<!�A�Wr����T�L�+1�$����;�c) �ʓ��,�8SzH$Li��{[7�y�	���P<+����t~B+�� �=�?v��Hҩ�Vj:|�YX�i9����f��<Y�#���8zU���-AQ&��Gl֟s�Z�n��8���῿�?���{JL��'������T�$�̾��A�j]#uL;C|��ݞ6`�C�w!<P�*��N �\a6���g�?ㆢ��탘Ф�b�������ȸ���۾ǒ�)?	�S$�v�;������~���	�tP�����5�N�"�����K�fj�T���X���]�x@����_qޏ2�ޯ}�&��a��o�
#��.2}J]�|����X0~i9��ca������ԙ��8��M@�0�뼒�N�,˿�E1:Æ�Y����&`ǽ(D��<U3�hF�/r�γ:��_qX����	"N�j���7��W�3ƹ�c��ý�	!qy����5!���YdU7���U�F:Q#0f���C�I"G��є�m
������9 ��-Bt����
���������n����@������}�v�9�u�J�.�$�TNp\���
��w�~��Wȭ�ro���9MPjFˢV���Ԋ��ufz͊6������S2�r�@�ᢧ��e���� �y�ںN��0��+�d��~�P���A������OI�Ͻ�  �pR��qOpϏ'd�����c#!�3�y��nD4�e>c�ۀc`��","��02�����#E�Σ���(�Kw8���Tv�"�-����={e��]k�z�Iwu!4/���Q�k�ټl\j��T�O`�:�C�}����#s��C���\���jxz���p�%&����/�����;���6^A���7L���J��(�_UWv�˽�4�	���Om����,Čp�L'r�����@�4�x��Q("vʸ*}ґsn�8W���Kմ�R�K�7g�8��g8��fwh�]h�T/@��G��G0��&�LQ�Ҥ[*�.<�p�7XQ���'��?�"5��>s����~w͉�2���W&�
"^�n7�V+��d%ΐ���4��j�Uq�����(�����4�xO(���3뵀g�n��\�>���g�U�ܻD�(��#Q�l.�+&�����ig
�9S.?�3e������K���@q�0��D�บ���*���3�43}5�_�iM����&C�jzkB��J*���I'n=�۹U>�x<[|�V&;͑%�`��O%�(_~&���x,��j��ۗ��K�rb3sY�J�������U�_�|ӝS�6�\��gj�Oۍ�s)޿���;���5�s8_�ב�&t��l��s�Y����D��?(�3I�4������y���f�1@��8��A��G�%ʶf^B�A��hB
���`IaB���2uo�{�?�w���+��3/Bċ�̈_���ټ����Fu�\�"]��53�OgXI�H������Ap���ɦү��#�$m�LB�K1h{r�-ʷ�����B�ΜPŒ�����X��dCs�>�\���k�"D���Ya���fu;�(J�ܝ'�� �y���^��ܿ��*��ZzO''6�	�e5 Z<>����XP'6+��u���w_�d?rq)�
Uȉ�4<OW� ��V����t9�e�w~l럦�B��^7KY��gE�+c�y%���	Ƕ��Ii9���i/��X^�iؐՂ���|��.f�&�x�>ч ,@�rG 2�}��Y)�Keݜ-�C븴v(	X���	{