XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��'W����d"�>n0Z�/D�t)�0����'k|����7��{���b����9z�8�L
��F�N�;Y��&��RM��}��`����_�ǭ0���&*W�q�4 �� �4��f4��u@�Px�O��LN�n�x�u�>���'p��u+�S�0W��~�^rC�U�>���V������zD�I���_ќ�S�Η.�%!��:^�u�>_@ȝ|O?K��^dK��rY��X�6�t�GP2NJ���~�Jٜ@պ�"6�'��P�b��J�X|x���݊j�_PĬr����ɽ�I��T#����0�\�YK[�U���1���`�;<�<"�L�v�{ŭ��:*�~���V��?��B8{�ჟĘO+#��.T�~�L\[����"@Y.������Ft�JKV��O\���!�������&I.��kHn	��n	��Л����<'���>��`���W2��$�a}�6(��0�K0�Hؑp�l��`G�w�"`�J�9U��^1Is��m�H�˂u��D2ę��7�J�r-��d�v�4/Yњ�u��htE���JH�s0oI����q*�w�c�P�U�ک�������G���	��5�N.�&#��8��� �m���mŖ�X�{�r-G��>hOl��Nf2��G4�J��؟�0�pw��3N~����I�]����fL% r8������A�Ja��<i�<��k��[���D�7�w���4�@,��r�Ȧkc᲋���5_�XlxVHYEB    3042     c80&�(K*�g�WqGi#�WC�pD�U���"��߆�&�=p
A�6�ITxD&&i���Er����/*�o���uh�U_�����H��s9�����꒯n�o�?2�߬�a�l���4�d�?Al{-)f�n���li*���$si	x�ݼ�o��.n),m��������6�ܙ�)^tj����7�g��{��hXu�BO��P���ʣ���.��ߋ&���ݻ L�/ǻsjx��9�F�13�Y��WE��3q҄6�4\;y����${�i�2�O~�����I8w�^^߶\+雱`�7h���?����BN�������.�G���?�ߢC�99�
#(��u���
D��*�%�����E" �-�zH�2�ى���V��$�ɷ��Ԅ��X�3�,���=��-�ܑ���^�6��P����"`I-{9�z~�O ��ߛ�w�[8�O�D@5R�`(�T���t������f�a���43^�~!Lq��ʲ��K���4}O�>	_������p��EN6��Ɂ@�r����%b��-���� ыg;L�;-���æ��$���P�����8�����:�Y���2���i���C��^c���X!�[��Ԗ�(�{ɖ�y~{é��� �ѐ��b���*��mA��B����ٺ�m���7P�	�A8����N����1Zu����o:��,�n¿���+u����Za�8�'�+���ӱ	D��1�`5��,j�Ic�1�����Lk�U��,%ގ�k��.fZ�2�QL�ry�иX64?ٓ1�Vj3v[g-���M����u7!=�g��Z>��ٔ���8��7!�@!{|�JGr�o�ҧ�Y����Ix�
�|0����^���Ő����@x�}��1( ��\qE܈tX�|n�g�9�*|\	E�k�����9�j�Z�ʥ�#�D�h�u��lo��n��ωz;W"������.3=jcIk*&Xa_Fj��ђj+Jp�@�u	|j-�'�t$v@��(�!Ò�ㇺC ���)�x܁�j��?�y?�Ep�[2��m�Y�g5�ܪ��'&�m� �F^�;�Ѧ��:�[��QR]�3�n{��D��d���wh2��Z�9�@t��j%�FG��u�`|	�`rZ��L43J+砾og�[���eJY~+G���~���0��%��|S��ĄIJ~�
����3Ox��4�1�8�?}k�K��,�iX!J���!J.����~k+��0�n"����8����G�z�\����I��y5~a��94�p�$����{�S5�b(Q�
6L���e��Y(z�A�,�&��7w}�V�J=�S\����g�_��Ð5�S�2�)x?�Tl���U��B1<Ю*�J����$�
� �@8���xSխg��
�&���V`Q������͋�A�X�O7 �P!�2�. ����M9fP,��ڻ��W[(/R{�4��5�XM!�D+�n�W:0�x:�͕�4�<~�67�%O�Bpt��_���� �v�բ��E���Rf�Q��NԊ�>�1x0J�+0�x��%�_W]gAT��9�.V[�����qb�� T?*)a±���e����2�MM��ِ���:e�3يM�2'^&��H٣��8������FY�P�ǈujk����XV���;�bRY���D�ח�&�+�ċ�;#+�����l�_��t��[�v���&w'����醧s|N*�a����~ �i;˫>�oV�Q���\pf2�f��4����(%����6p�;1F�J�#r�PITeY(��U��N��v�_���60O�A픠��ݚW�S+���B
��>�dæi9�����}d�7q����c9���.�$�s�Ś�����}�3�E�ǝ���N��c.�#���	4/�CL}�ɇ����FUo����v&��F<4.j:�bK�B�l�o#F�t����I �M�zl.-��W@�g�^݁�~]
�ȳ��6<C`OI�~�X~�э� �Xg��+Uh4@�J�����o5���+W��d�t%ݷo������L=��}�~]�9+����7.=�0�t%�.ŏ�S���R�#4��ܨ�'88�s^����XmE���!��~��p)�=����4��0.=���͉R�N�:giW8e2b��l�� �YψA_�s/�$��I���Ӛ�'4m�oT���/�D��@*d�-�R�Mv?7�§K/����I���N�%'`7�����ܮ6t7�! �o����l�� ���j)�
���� ���M�&������A���8K,+�|���x�@fBN����C2C䫑��� ��^(��	R�O����lb�qWSf1�`�!��۟�#�΀�����g^�V�_�K��KƑ.��"{ǿ�͵|3E5��,�����l��S2�(	���d���{ˤ-1�#f3�&$]z�j���H�m�h�UQ3箘�,)�C��JK���n��r.hI/�E�^V&P�đ)�l��Q�M����Wgޔ����}��[���]JQ������=�m]�	h>���q���S���W���)l����9Kea^ȍ����x�0�0L1�0dx"�G�7L8����	���h��)V�b��𳩨/���T��l7��C���))Uܤ�A�
~Zom�Lb��v!��I`�7.x������jц��,�Yx�CѣT�ܻi����\�C�~�V�X�D{�>����d���.��ó�X%�Sm�5*+v�o�vn�L;��\���!x*2��M�?J�O����=��7���=wd�3Sh����iwR�
[G�ŭz��%�,`�f�k~�I1��l/���'}d�A�c���Y�&w�UI:�8Ug3�������2��9m]N)s�&���N�4���6![��>��ے{6Ə����k��{*x�g*%�}U��i{5$�*�^Ve��׈�-;} �]zΣ42�;tH~�ug,�
;�t�&���b�8lm�õ� ��p��m��}��'�`f_��&|Qxhp<.�����ffP�P�j5�\a�B�QW%\���-�ߺ�)�Y��Ӥ��}�b$��p#��o�Q'W