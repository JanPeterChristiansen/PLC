XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��	t��:X�U�����v�A�;Ĝ\�\�����`��0�^E�KJG9�&<��k+�Knݽ�����Kc������=�N�<"�=ɏ���ϩ���g�S�-j�o��wlo>�8�"Fw9��b���n}�l�FI��#s�)�[��ީ :��W��%��vmR��Q���vl�<�kX�Z%�NN�mH�yg	-T��P'�u�I�˞���B;��Յ�2{�H� �]��%s'�R�����܅�E�8�ĝ�m/�R] ���u��9O1���e��^�c�_�,7�z]��LV�NA�����������L�Ne�l*�d���-& �RPF��c�~�w&Wꖊc�x��֐�H1\=���>�@�x��r�8C?�6
�>�0-��\KW(6 4֐��ĳ�f�[,7��0�qNW�`J�J5��?f�*_fB���?Ԁ��h-��u�}�͸��1n�;�ǝ����
���wz;���5Ȭ�E�e��e���O6�Y��Z}j!Q_���;�Z�O��+��,��g���]e�eY�X F�xa�g6��!Y�Щb�*���e��r��?:��[9m�L�������(ƪ#`�>�2$WVVU�d�/v ��W�R`��h�������љ�#-PW��|�F�Ѳj?!3�`���!��D��� f����>��|�ձ���H���~D]�[>5[�_���

܎w!�#��xق���cw{:�nL��!~̾�faN�Kٮ���*ᒢ崙�������Oj�� �vXlxVHYEB    fa00    20305a���-�CQ%�q��Sg��d��ji�'s�;�p�O�1�[ILuvW%���G|�T1~`<(��A��E��%�+�`M*g:J�Y��oѿ(���
�3��3D�xDh7>6�G���ӭK'�~?6���F��Z��\��P�G��{�5�a1f��[�=�ը���w�\��]h�;Z-�)�o�f�2'b��v^vI��:p'�PCU����zf�����d��l��&� ;�XD�[�u�o���nyUص�Zjx+�1�ؐ���� |N�)�V+��+�M@B��x8�5m�ƏH�����Y�d�w�QiX��O)[!7;x��Q����y�|��ի�>gc#�Y�����2h��n{%wS�$���9`|�ٔ��5��2<YjqO�()xnJ�n�K�O8�3/ ��s���'3���B��<�:+~ �?�h�B��Ӣ6�En��Aϖ���sܭ3���|Q�?`2�0�%ws0��=�Ӓ��\.3�{
��&4���
�BT���!�.9o�I'j����q��F���Zf?d;u��CXH]��d1�!���z�u���ZL�g��޹�ʙ��Heo���l��h�$b0�8�-�jf����ц�T����޵
��%��U�re]��G��������g%JR�f����1Ax7Җ�s@�ƍ ���E�mU"(!+|�\�ǩ��Z��)����F���f��q!&�f����L�\�����y�_�B�С��}A9X����b�Y�$ؒ��H����Y��,Ԋ�&�#��R3`8=Ť	����J�p����8d�<";
jZE��5�&(���#m�� m"��UA��x2�)�'�o�]y=��[��t��\�����%Pud�\������T��$s��B��D�\�)�_�=U�簲�ࡐD��q(�b@ƌ�i�����/Ee�xeN�u�p�}��D��3����� �?@��l�U�F�F:��l*��m��63����H��gAs|r�<oG���G镯l� ��Cg�U(7^b����>�ӫE����y%�aT�a�M�C�Ԛ�4�@X�uݳK^�������G �VCqU)�����hK�=K�5XW���4��芀F��)�3ӵ{�B�1�9�*��#9(X7����['�*y�S9KfB�|�b�h>�apd����`��\fK��f�Z��h�"ě[�����*C�^��,omyP��v��޳1 ���j�<�z:� X8�܄?��C)(1����w���57L���n����l��x(r#�޴�*���������'�*E�k�A���'�j?����]�7�q�X<t>�6+8�S�������4<�t�35n��Bc`/`tx��!�I|+�r����$S��F�)K)(eO�q=m'����N�8�{]�7�a ����O��Ǝ�,W�3�̩��N?��%H/�7�S���ޫ\(�Xyo5�g�_�3atj�<��^����V逿�jj�Kzt�o��T[O	n�4���6H��� g��i�`��ݵe�d��I��M������q�<���{�q=@��(�9]5��-��u'zjf\$�,�{;�q��yG��s�� =zh�D4$���UVv�<�MRe-l_�G��t<%=htLm3���4�+�\ە98	z<&�S\n���xT
��;m���c&���������B�2x~���ؐc� �j��b�����1dG���h�'���Y]ZdhL�k�:���u���?��k��pw��-�p��y`���lY<���Z3��^���[�T��*1u?x�T.y���δr0�	��#�9}��=+��~�5���
ɰ](�j�?��#�^Z}���Աx@O͂9|�ˊW6 
�`��=��`�VNk���?e�Ɗ[~�O`���K���w����.��d2z�m,t���W.�R���?gs�kP�y�d�����╔Q�!F�j'�'�޻��e�?�r�M@�n��&�HR/GB���
��1�o������ll�$ �͜d�=X�� $��s������T����A�m�
|�R�����b�I�}�3*c���$��8�-��n2 ��$Ǻ��q���Z$N�#�j����~�(��I�0�_�Č�z�F]W�׆*vn�FT�mڡ�}����kG��fզ�<d��M����n��3'2pG��ߗ���r������]�Z�)����q�ȑ���;'�i������Ǡ�>6f���M�B��,����R0<1�a6�ބoC�|]�kY�p��jF� gI7N}{�Q����pc<w�]Xz�ڨ��g�n�Ff���3駵��@�����Y���Mb ��aH1�'q�?=��,9{�P�N���w)��>*%��>eK�l���[ĝz/��v����ɐ�����?^��]��L��vݱ�;7`��/_�6z�;�^�{	��2'�f��+!'�^}�������� ;.��:��bU�1�z��ЈU�T%�W��
��h��Xy`��������%n���IU	��.m��x�y����EU�)����r��lk�f��GI"�ʁ��B���Aax��=�z�����n,_�j�<�t�33zL.+V�]�����G>^��yKS��]�C�,�p��QM�5-���u��rt���4�Ç]�t����[P0t���Scﯻ�����bf��L%WE�h[�c��γ�8�XU�H�Yܜ�@���*1B��DDMa��rğ\�FP��Nʋp;�/?<�&g:��K��l-(k8c��s�in��#ۥL�r�-X^<�M�8Έ����C�Eғ� -H�Hyc�h���_����������)�H ۸)۹�on��{�w�젾(����f]������
_1-u����eϑs�fML�L��/0����p�)W��܌(�ݪ4����m���2؇�����kJ��ؗ�Z�Yb������2jX%/�d�T"�25�����Y2)UI�50�~AN����˾���2k�;-R>���HY��������3D�79)E���3:TE��M]�ڐ�/�9��T|d~^�#(�S����Mb����'@�f�kMh��Ґ�٭�.k�߼�v��ӏ&ż#}6����"@_R�]�'��s�f������O���]��Z��M���hǷ
�H���H �����cq%��8y$_�D�ShU
&-�6w�YR.m���I*��&��Y>	�<��3�b���h[���[zؒ��3ƾP�˰�ߙ���׆`��Eڻ{�F�hh!t����c!�Sj�`��>�x&�!�����լ�~��,�B&V�a��H��K�N����&���oU�(	:�?r����t��*s�G�?����&u�f�9�G���y����'��M���T&�B�gB���%7���;�Q@��;oP��LF��p�a>!����Z��\�4sLy�v���Dە7��x�ޕ��J�(?Z�Iȣ���(M�����\ⴔ��Z^Ϯ�H.�j%�j�:嗱��������KyC@���<�腴�t�A,��6�V�AP,ٹ>|���>�_fI�Z5��=����n���Of��\����:!��r���6�I���,�8�,&<)1�8W`j����F�.^w I��
R��D�Ո|d��P6�(���a�4&Ie�4u�i��7��?�_�L�&�xNvp�m�H�ߚf�7B>�ϥN�n�ο:i+��s�v����3�]꟢�c��llCiS3�W��ᴕ����*��m��xR�OE��Os}	�%p���� i2�i����yL��O���+����W�a{��R��]�aEϪ�����7�<���3��B�� �|dj�U�*��K��_v㟧j8�u�)p�`|�׶d���ܵz2ԮUE��V����8��R�����/��9H�7�t�	��I�f.��<D�/т��A%��0{"tǠ��{�������X�,!��)+�e��3���I��l	�O>������.�7;@���05�r��s��&�wQ'�Ŕ+ɽ�+]lA�%[�ɋ���|��XDd�"�f=t@�V��4��L�ݺsM4�Z���/�;�"Z�S��ԁW�a8��4F�0aE_)���eYw��X�L�>7�������̨7��cQ�}ߑ@EѶ�� �.��D��������W�n2h�*e�~u�SQ��@h�/Dje�=5��2˭zzy=g�o]\��Z�"�8�2���-H�1�����u8��n#av~����'�|�l���O�W:�"�(QQ���]��w-!:n�b���>�������Yf�J��7��⦏	���L��剆ˁ�5���A��!eLGS�J�)��DZԎj���w�yYV�0aм��\�/�|j -뛅�)��흾n�q�Ee�AVy�z�5E�e�%S���|$)�Cz�xg��h���<HЈl��m"1O.l�.�z�� ������d��fo��yjA��,�N��ӄP�j^�qI4���f�g��91�Zc��9��vҠ��Y~>D�c�?#�/��X���W��Wp~V���pPG���&g���C �~����,��-WX�ލ�1^a}�f1`JJ~��1�xfFg:W�K��ն��´8B����*��=�τ`V�>�.�Jz���A�\�љ�V�*��|��Y&���F��;����3��-���q��g;�Q�{:'8���+Cr�;F{'߼�0�û���|u��3���_Q�6��m����IoPM��,L�c�ב�f �s�f�\ci�����������S�P�ĥ�l�����Ȱ�؈p_����ͧh�W��~�����y7�h��Q����kb�Q�BU=�"��bՎ�%d�QU[�/�Z�.ոv�QF�X�1� Jsz�mB�&.�T���Z&>�d�![�����P�1 c����xtcw��+�,{Ϧ�Ԥ�-#%�m��y��u�"賰���8��>W��U��3D�r�5s��{�Q�w�WRT�J*��,M�,�e*��Q"D�rȼb�R�jE�������JkPw�c�x����/�rdD��;D���V��.z���a�[ő�ׯ��khŝ�<�@���]DQ��4Ǥw;<_�ɻO��96=̔u�yE?�`���Ǳb+#�}����cX��22o�$���>W��PX���SGx7UW"�̉%R�����f��&y�\ԹϚ7!����ѝ��K�dC� o�{Bg \qQ�3( �>��R��#��b���<�#�JKĿR��9���`;�8#�`==�B�����s�_9���=*�l���g�zJ�dY��kn�����]�����=՚6�a����|鿰�B�If�v�_��zB2��5�W�E���n�S;�ZR���QR�x��m�B_��@U��	m� 7�!]�MS����_�H|��
�� �?E�w*��`M��z¦:L���庸�!+�Vy9_e5�<�����!�Tps�9ʋ��x��
9����C0���ȉ͈���YQ��c�}���֫��0�n
���id�OK���&�w��[���N�q�3h���yл2�����Y��,Q�qr4�J�g��8*�o�t �KšY��N������W%�V^S=�H��j��x�g������bR*�۠�UL�r�<�6&�mՍK�y&R;?[q��S����7e|Y�܆ć˃g�����~��N��W-*� �5u_�D�z����rĕ?ԳD��w�?C�t��OM�c��R9W����l�����y�^)���qɪB�"�<l*8���i�s����	6 gȴ?�I`�-�c)����W�GDXJ�-g��'1q8�b��2��]����ߗP�e���`�V��*]ܡP�΁�B�����?�"S���Qо�H'��;.�\�����ߌ̷�N�i��q$f�Q����s����#����@|��:7�u\�b�����;�-���l�dd�'B�Q����+�o�jTF�0�ݭ����������{�d�n���>I��gĵ�_�dP�%���:*8��8E���1j6�p��(z��}i%�g%�r�g��=�z@���m�j�Xw�2�EZ�{�=҅ȲO�D�CE^43#���Xֲ���C�=<9��O�c�rm ��=���5K�5�|9xf�qL-���܏-�	��Ph�N�G
\�Ҡ=�~B��T!Č~��N�&n�3�r6u��I�G�������{���v�%�7h�ˠ���}V���X��a�?�꟨�!���cBm���
#��R� ]&�0[㺘�+��3ܙXaM�1hc^��ץ[n��s��/�-]�ԋ�/rB�`~��7�WD+�&�s�L�ְN	]��}/����,[�d�
1K:���D��w�Ή�CZ����n�.:�/�W������M��^�w��\x)?Y(������h^����N��������#g��.^{X�pK���8����x���8D�����؂�O��+K"�����K���F�����>��,���������3��:�Ǥ{N�ޜ]-SZZ�߱|�um1�iZ]cc?AYUM�2���2FL�A��Y��nA��D	���b��H��YOZ�Q׏����t���.-�]t����T�d�����Q=���{K}����C�7��j![hka�Nf
7�
��s�}{D����>��Z\��(u�E��o!�,�z �*z������͟�I��*�ę��p=���=R�5�q_B-����=��_����ut�֚š�W�V�&;�,�M�	$�-q�
�0�ˆ��[��F^?�(���#M�q����i/Y�'���ϳ����H����p7�g�����۠3�اR�vc��hN�D.��e	��1�D��̌Y��l�y��zk�u��Ɏ\�G1*�̳x�8��`���0y����'Z5Цy���MɴZ����ᡛE$n��.�ȣ�3�">�vd3>Rg/ƿ:�fU�lYu�٩0��������Zߴ��W��<�������wy�	R�/��z���&����0@���|)˩/o�}ڲA�L��`���.r��y�jޜD^&���b�b6�?�'(]c	Q`�66�_i,�gyl��}]qY�aa��$�g�Y��]��������=����F��NI@X�8 Xd�I#�Ӫ����臘��*��E�a̱����i*Z=�a�|��k�vP0�z���f�3�G�Z2fJO�� �Mll^��9qDf\mN�P��*�B�V�Q�0�󘣠�G��B1�eԽb7��_ʽ�!1z'�n������	H�,c[-L�2��|��hg��$��}���}o6"�����t͒%Z�쯱���ۜ� �~,��:�
���KuSS�����Hu]_�P�J����fI5_�o��Lhy9Nc$�F3E�Ĺ��Q4A�i���W���\����O�I�l�Ě�m+F�ٶ�𗩠��b)�p��ʕbN1as�B��(`�ŋ�ފ�2Cc�[o���0�ͱ�R^SxF�"N�0�s�{��܌�qo���^T��ր��X������!�uy6eۦȧ��Mݖ=)�fa������)>ս��5l�niR?+>K	��R������|I��M�h\Ww�A+�%�8��4�����s�=��(�1(����~��M募�:vI��Lㅞ�+����wd�;����)F2�
�"�h���Δ�����jG�Ǻ�,�{v�±�Aj���}*p5�d&�˃]o���(L5������Z< G��K����i)��R1S� ��rfj;u��fP9]p���v�<4�Qu4Cȿ����+�>D����X���*��Z����p��00����I[wܸ��` �DC'0�xO�����^���֑����.r�(���-���3};5?����u#s �R�)���C��T��|�v�&%����s(�u��r<H~OᎪP��WW�ad�MIb��6�ι^���2ĳ|6��]��B]��ت�H�)*r���Rk�q����'���M}#jD��7v!����M�l����'4!}X{ѐ�q9��j��եO+1'm�����N�FXlxVHYEB    9620     d70��/��{@�ݯ��֢�u��i��X\s?Uey�ƽ�?T	{q�>�D��(t�)F����gn��ޭ��lq���r��S�\Dɤ������K�ó����h#��Җ���B[��˪!WU�ۯ��ܲ�ח���� ���Z����������4����X��<ǙvmrT2j���)�h�?�v*`֊'����BA��+���|�6�Qmj����M�#Z���;|�%M��?Rw�DF�n:6�_��u��#�H �ƾ%��!��]K]����2"r��E�Ʌ�}��1�
5���}��ב 9����e�6x<Lw._����:1��V��[�����p����~�:�W�%��|��d)���%��������\
�>�FUhX���R��UD�dlԊ4Q,�ً&<L8a���H��<��q1�;_s}�&x�ܓg	� 1����5�sh?Y��e	ìPGp�� >x!���O��
Ӧ��.t�%i�z�f��g��w�I�<�h\1�����$��rc�LYh����)n
�K깪��#��}�^t%�7���ڶU�-K�Oz,q�p4��,���T��&��(�y��P�_�ʱ�G�d�ۧM�ae��������M&,�[듴<���7A�j-P3Z��Dd7f[Q?�j�4�-�H��nu}�f'.:)�@��勔�lZ��l'��;�v������u����0{�6g!��X<�jd6.K*h�}��������ANQg�����;���z�[�b��
�%3eD0؟�&�T>X%�9)	��/ꀨ9I��6�Z̐���� 5ix Գk��&�n��T�B_�F��`�n� �q�(���jƦb���8�F�1זZ��f�{o�֟j�B`��?�ڲ?G�@a���.�ԔF������Jm��MJ4%`���:ͯs� 㜯�]���{�����C�Kh׉q�U�=|���l̓e�$�6���>$��ȴ�����;�� %�FV��]A�mjB�qR��8]P�3z��]r�����DR}�5���� �_}I�`�	�"��BVt�#���
@o�����r��?l�c �}�\�:�ЦӼ'�6�����k��hV��ȴΐ6 =��eUʸ
*j�x���W��NW2x�A$I�묁���|�~r0k�X'fU��{W���%�r������a���;���G/gh�%�sΦ�#�߫ W�:�po�,��g�����0֑
���<�gW�:1X�{㇞d�a��se"E�Q����RPM�xĚ,��z;�{�Xx'��Ls�^VŰ�:հR����^�ȷ����-���O��L������LBiB#t�����嗨?䌝�������ǚZ�  �#�V���b\�;!DST���\?������Tbn��ȝ
��P�*��?*��nd���&>�_|�@��L��dݎ0��'5C���*�Хv��8�Ux�eco&\z�Q�<!��k�\ďx�5�חn�
��AS�3,���2�G?�ĸ����,y�8Zx�Y�y8	�a�B��\�)��绖r�/�1���_=?^:R|L��z^x<�:���к ��h,[��1���DI��)�\!�R��/�W�J�A�&E�s��QXM�n��W����hbe
�����η��۫5�5��K���,��O�#;�I�bkz4��ң�5r�b�=��vщS�@�U�?7[�6��|��p�Q��,��5�5�j�L ��[TR�`��'Ƨᵓ�,�!�@?�_p��y�z�xH�\��VI�q����JG���n���y�Φa�w;��9`⿉�|�F��f�Ӛu������*�Ta9��.'Y
���}R����on���(�J�ɪVT�u{�Y�
aǏZ�6%�0+gb����i���b.�|��2���?mmp�j�Nb��m���	v tL�������י�)0���,��owv
K�}y�6�x4.�)mH*��������"��l����t�w�b�'��o�W|��j}�yv$��.��i�+�</���)�u_c�d˜:P�*�N���n'��GTϕ��O>X�8�Qs?�����4p��_M9����1�Pŷ�ULa��z;V1?Z��@b����5ʣ*�t�T��a5.���}��{<�PR�7��\�S�����9�f��?��!�>��0��:�2��{�(�>3z�I(��M����T������<��^ׂ�l�}����)�#+S�y`����᳥��<����w1!A�~>X������M��C�f�ʦ��J�){s/�͹�"���ۙ粲��4j[��kwd�%P�X����ƹ ������K\��%��2���n���4#�����`<z�����h!Z2�7�Gա$XalB�:�e2�!�ǌ�_ε(i�5^ztB�~�1�J{�`>����+5RBrTe�ȱ���6'��/f��n���;vpI�~E��Y%;!��t��(kH�qE�R)A͚m���_�<ϡ*��2������ȓ�:�?�(#]_̲q�8%P��ƽ2[^�m9>�!8��=���$P�/��pÝ�u�4(���;���+�!���#�%�Y殆ũʦ���=��WS^���'��y �0�B����~4Dh�$t�@��⧗~�$Zu��_���;U�W|�ҳ���H~b���Ͼ>擩���ŉ�ܯ�2h�y�:��Pu�շ�����ջy�bK��@Ei�o&��j��b˩X�%�K���K_J�~��<&�^�=4�}#�a�H��	/~�G�X�Y�!�����N7^�/�9��^-��݁������$Q� n��#S.u�=�D3��գф�$c��g*;sʟ7���q��"^�ĵ.������PJ'�Lk�_څ�ۚ^W�q�r��q�x�ǘ?ޥ�1�����Rm6���t�'�ﺕ_�M:�_m�_�5łz�_\�1T����B�mV�W�0��1��^9,<_h[*oȮ�� �*x�����W3���y j�8ic������(����*Zhk�.Jc��bRЙ#%dQm�L���}ǳ\΄�?Z�T�^4~�%!qCߴg�E7���]�햜X+{�9r�G����B(�t��9��36�������_�`��/����P����m��ݍ꿶D��e��L��E�Ȑ���
0ɏO�@��ӛ\�03֚
$/~fp0E�ӑ�[c��B/�):KW*���Q��pL�NYBi�����F�������ѐ�)�;�0��7���DM���t�Z��F�aQ�,0@$����+4�%���q��޼B���b�iƖ>d~�;$U[��Z 7&�Ϛ�A/�