XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������:0�O�����ܥ��x�y8��9����;r�c>���-��_U�VY�Ӫ}f{[9��B��W�`<]��䥤�:�����@��B#�.t,�� �'��?�x��J�	����L_�T���Ѽ˯E@���Xq��t��z@O��+|���q�c�ŉ���/�'�2ώ�Zo>�ٛ�X��ع�w�0j;=ɺ�~hF ��7�)4�~��e�s�=y�P�du�u��0���:�e��|E�H>A�U�~�[z�ؽ/k���ێ|nO��p�)f���MW���dC��6L
���C<{cv�h�u1�FX*��8����Z�ҝ3�d��p!�c��v����0�(ڳ�ߞ�ȃ���(����ҝp�En�_r�~���0)#�̹��#�E��k(*3��{�E���wd;�'y��R�����1�:�[�[*K:�;�Q4�y��uz-@��S���6'�~�
 Y漂�˅�'B����t�G��x�����*�qH����d����~s�٫#�ۥ�"u�4�2&2n�uV��s���t��К�g���XD6V	���)�䇄�=�,��CT#���3�o���[G\��n�:I�w�~�I���hyk�RV��9]���<���Ʒ�Rx�Y��";�3���=���ႚ���i؝O�Q��9�}�X�rt��@!�w�=�ɱC}ڤc�eq�Cb? %�{�	i����GU�u=��؞�B��Qx����=3~����?�5�5�z)'!����yyƝ�XlxVHYEB    162c     850n���ߊ{k�o1��τ��-_��׈���l�a����jIJ��JRX�!^u�?[�^x�AǴ�5�D����a�F4��k�E��,B�#�X�Y^D��쫞a�_�v4z
�Y��1�Kn�4�F��ꌧWv(W��(�������1a�Y!���i%�]��]���f���-v�z
E#�d���<��@���g/�\��+�v���\n�'5.����9@7����5L�a{��m8��@�e�z��b�f��@�ȐEq��u����Ӂv�8��s�@}7NNV4���t��x7wF������Xv�rbp0]b&T���\����}�W��>���4��լ�o��)p�n�8�"���5]��(��>���b����$� �'�U5 7"k=�$*SB4����ʽM<����/d?���V6���M�"�#�H�]��x=�������4b�k�����<���kӾ���2�xF�|�o��k<cVp��aC�:�O�:߯<���jr-����sh�Cx�����*�� u�S���J5��-+Ї/5��Ft�� >�t�̦��sB��c��Do����o�����۫�p�����4R��xTd�����mh`�<r�{�@��K�%.w��(���g��Ry��柋�Ic�H�C^�k�ݘy�1x������a_���$�ü�f��^����]��Z~W�4���ZD�wq���pd�Zj�u�'�������mr#������6�0�8�a�%�����Eb&�����K����ƽF`��C����� q�9^��y�(�x�[@O�ww�պR�*7l�?蠆�C�����iэ����Sq�I���>=ιt�0�K���-kL����яԮ�q�Տ�DM�Xu��|�����Ĵ�qRvT����T��s����	�Q��(��s(�0HnM�y�6�zs��y����-��B��Q��&��qa����ۃ|1�i�1"ډ���5Q.݁�[���3y��|3˓$v�~ؔ�\����G��`Q��UreL �����G���FG̝\�z�݃�g{��?�ZsC�����N32nQ�>ؾ���#��[M�d�ן��)��a���L�z���TkLe/����� �۞#�·iA$@b$i;l��e�P^
2!J�����ͣU@Tv9h�D�v"�N&�7��@!�3}�8��3��^m��r�IG@�s:�C
�I8!{؜�_���j�]nVsden��݉W_ulUG��ьV��u:n����{�ϿI�1]/-z�$r��.��F�F�{�R%s�>#����l�E��UN?�?���	h<���U^��]f��9�������:������i&�Ȏy�\�=�a��ե����uG_��^�<W��9BHV�Tdy���s�x���\�i垃S�S�^EE�?��閊�:m<�����MG5�������Օ5�+_}5;+qEl(�܄��v�!�)�>��0�5���f\������Ǩ˧ؓ��<��v!P��s���߲�<H�Lw���6k���],An�}(��ƹ k?��l
'�+�D��ٹ4������=���9�U�� 9��c��:E"OO�j�����h�
 �F*z['�?�8zT��]{�.`2\ߴ�f��Fu������<��p�|��A?�|�l�'e*�saF�	R����[`����O%���) �)����^
ސ����05f�Cf��v���H�]ѱ���Kk��� p+�6�&d�t\�P>�Ĩ�f������'�2kh��F#�j��{e�*v�g[}N}������i�e�$��o:�+ث^q��9î�i	3�wf���_�%ŹP�u�u�7�����J���{>-�Ը�'A(���\�l��\�"��U�4,�L{c��v���m꒟^ѝe���o�փ�?�uz����V���7�JX�r{�n�@/� ��$�͆�֌2�3ȿ�u�}�h�l/e�,�Y?w�_��Շ ��G����O<����wuϪ@^)�C���̗&����TG�}#�;"��*xEz�k����F%���w�� �_
Չ�jx K폘M��n�#h{�Ҹ�