XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��B��B(�u�QU�Q��Y�ˮ�j܄��,��{{Ԅ�P�a�Lu�;��
�)�V�.���=��:�ӽ]8I���J!:V{��F��mc�a���'���c������,�j�Z'Z���Nkb���x��2�AW�X��R�v��OD%����c��V�S@�3�C�M�]@V�-I�~��{U<���z��n�hCS��h�����8_������f���U)��˨A�	X!��4��u�S�h�&�Q���P��*�ε'J{�}=s�[%I���F�� )�1�vO>*e�k�e��o!~���Vʌ��I���=��[����<e��H�Al�7z��c��a���r��N���+���t�Ǎ!�ȸ��U(R�|�#
+��\sE2�������r��}�zuT��ݢf+ĴCU��[C�5	;'ִ�D����H������ѣ�﫸A Έ>Q/�lY�� �	� A��>�X��L#��Iw� �������fY�>��_��F"�U�.���ӻvO�P0���	lW<\�*R��8A�w�l�%|����k��h��$s9#[7�_�~$m�wX?g��F.6��Rb��Nc�1B��@�ec9a�2mb��6CF^Uq�/�q��Ǔ���r�iy�r5,F�X�����H2��+�ʜ��Qt?�tw���"1��R��@!�<�/5Y��`�?�7c�?5_����g�m�'�0Ss�����h��LFJ�*W�gGJ�X� ���rZ͓��7�г�
o�&E>��/Zh�s�eİݖ�XlxVHYEB    3504     cb0�䑿4}"D�bB"&fQv�Ah��Wf��*]����l�jc��O��z���Fl�L6��f�jʡn�CZ��Fh3��:��biX`��)�ޞ0�jU��a�� �/�a���la-I�V�D׍���>3(d|�0�������2�5bw���|ȗ|(^�b+�V.���"��I䵦j��=o�h�vfn��x��޽+|�XO�۶Z�{kn0��g&{u��\t!+Q,2&4J�78t��B�*���)�9	8zBJ�l�U)��"�KY��v�@��' u��� bPs1L5?�'�"~O�~)s�&��2��!>�'y��EP2��0�����U�S#O�-&@��SF��_��j2=���	��6�d�#�!�ョǡ�\{�P6����-3Ni ���OV��>�@ε�_�6�H�g��+BC+�\�Ć%x�|3:������� ]�h.���V�r��V^f��&�H��sB��d�̺���b�C�x���W���ɠ��*KR�N����&���x��_������]�/����徹a�\���BGE�Kg�����OV*�]޴�ѿz}��F˝]��:b�U�u4��G��x*�j@z��bH[O�94zd��o�f[bR�E����<���h�❚x��S�x���Hz��rB��� ٣+�{~Z�Ck���K�::�gI!~W�-�c�����t%6J�ᶼѺ�꩹0�#�:*���E����IЪ"F�%���
ߌ�Gl�?�#pP�>��i��`�V�X�_��9��1�ռq��6��S�{��r&vD缰vmtL��®�ǻlު����]&(ts�qp��L�ܟ�`��������8d�%������+">��Vf�$&^�Z��UYz+pM�d�n�?�n\������(Q�;Og�Y"�l��C�K��m}D�5=(PU�mI5����/ol��N�T�&񮹼�i���$7&�	��N�5S!R)�]r�5\_2�r����u����VC��ݾ1��n�pf}�̤̐I�"J�����,b�!eԤ>F�l�j��uwƯw��)�:@I�x����-YB�>�q&�bű��G�&��+,� $l�T��9&����ˢU��o�OZ����uz� 4�kP����<E���#�6���q^��lJ����aD�id��|%*������Y-|g��սd���l˩c�v���jn���G�fC�vGTb�Kf;W[�P*��ڰ;Կ���<f�kQ�ɛ��r@�6'S�koل�N�dC/뼢��#�i�\>Ǜ,_}�*��Ժr�e�	A�|���݃��[�>��%���n!g{��� �`(��o9��S�}RR��" �!��tya��2ǒ�\��}!�9@�!����g�?�|s� �j����S솿��a9���J �U�@�=��2�n\_,��;�u�v�m��/�,�(kٺ�˶p	yC�&"[�l��3խ8�j�Q���~!
��.vSP�n�� 1�S��l6^�����\��G��r�K^8V����iW!�K�?ԑ4����$ǹ�O�H�X
R�0���ym�.x�Ms��|����O^�ci�"!,RO��-��8��F<U�8�T"y�6��vC2aؙ�5��&�W�c\'�D���m�Ԡ�$@�{*G��2�*���9��?��8�������8b�� �(��ʻ�ǰ�ޡ'[����u�����?2��'.�"׋e��cT�ݍ���ha|z����X���<��ڍfUe�'������!ݸ���©5�_�����x8���.�N�IX���w�ȡ,��|<�-�R>!YoL����N�f��1�5���t���~F=V�v��Ϫ�m�b4ģ���M�z�����������KLa�ʣ�zy[�N���^�8Q�Oܷ��N#�7cmT��|��n��lU�u8͵�� [/l�W��pF��v��O�I]�(��ַH[-�������շL�����������΢{	#Ok3)��FO3k�`��3��ŁE�a���U�0;A���c�����Y^�RMVq�:����tݼ@g{�~�8�W��E����}�D��'?v������2�:�o��Z����I�g�e�P'�dzڄ .j;���E�WO�9�?�Kvu�ȷ�,�����s��Y�tB2��\OĿ��{i�����K9=����|� �J8^Tfʏ����.4�Z�n�!�P�v�4�.�F݃��w_>j[�~\R��g��w�g�u8�؁M�n�����;���k�rU�	�#�1[����6�6��F �U�� �Z����n(��T%�,�RQ*wn0�O���*?�S�/$3�n���֩�"��P+��t���`ol�O}�i�횞D�8��5��*Қ8j���2+����M'��&�G��4�o0փ���'��c����^���ʿ�	:1�'pؤ5::_�{���.~�+���<�8�ݗL���|�7�qڤ}1�tճF'~$�?��>����?�u73[����e����6����WՉ''�=V��-8_)�¬��ePǛ��M���D �bͷA�&�����%����G�!��?#��+�Wo�`H\L�i1:���������t�[��M�%���w�_���`�"�n��O���Bʴ!H=�	SK�;�Ϧϰ�@�<����Gf��ӷM�3�p�&�t�}��n,��N��Q�!�9��l�AMK�Ȯ0r]�� l�&5/+�U��p/�6��m)1{0/W���8�LW�=�Dﵕ��@�u�g��P�810�L		A�b�+�W��|��_!�X��H]7-_V�� B�5���Y(���*���Wpw<]�����L6��[�&3�e�m����5ex��SUQU)UF�z^F�f$!Ն墤{<aב��Lҷ�B�zS�{ ������~�Z�����䔒���ӡi�M�Ύ���j�����@?�=@���3Ż�`˞���
��rB���lL�r����?�g *j�h'�#�u���j��h�T��L�2(x�𖡫�E�3Կ�gL52[&E�I���"U$mFh�U��L�������u����z�/Š�ݤ����?�pU�$g��Q�m���86)���|\������(�0"�������V|8�ͷ�D~�3�$�?�J�[$$P^^/�Ѵ�Qu�/+�THV�م��i$�$��2��߃�6~5